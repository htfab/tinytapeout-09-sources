magic
tech sky130A
magscale 1 2
timestamp 1730795883
<< pwell >>
rect 3178 3440 3230 3492
<< locali >>
rect 2936 2440 3562 2490
rect 2936 2202 2984 2440
rect 2212 2052 2984 2202
rect 3508 2052 3562 2440
rect 2212 2014 3562 2052
rect 2936 2004 3562 2014
<< viali >>
rect 2984 2052 3508 2440
<< metal1 >>
rect 800 0 900 100 0
rect 1000 0 1100 100 0
rect -9600 13122 -8604 13310
rect -6604 13110 -5608 13298
rect -3582 13114 -2586 13302
rect -592 13122 404 13310
rect -11158 12894 -11152 12946
rect -11100 12894 -11094 12946
rect -8135 12901 -8129 12953
rect -8077 12901 -8071 12953
rect -5146 12900 -5140 12952
rect -5088 12900 -5082 12952
rect -2135 12903 -2129 12955
rect -2077 12903 -2071 12955
rect 2438 12714 3142 13306
rect 3074 12108 3142 12598
rect 3074 12084 3176 12108
rect 3074 12032 3100 12084
rect 3152 12032 3176 12084
rect 3074 12006 3176 12032
rect 3074 11518 3142 12006
rect -10470 11364 -10464 11416
rect -10412 11364 -10406 11416
rect -7428 11370 -7422 11422
rect -7370 11370 -7364 11422
rect -4440 11364 -4434 11416
rect -4382 11364 -4376 11416
rect -1440 11356 -1434 11408
rect -1382 11356 -1376 11408
rect 840 11390 846 11442
rect 898 11390 904 11442
rect 1546 11374 1552 11426
rect 1604 11374 1610 11426
rect 3074 10966 3144 11404
rect 3072 10884 3146 10966
rect 3072 10870 3182 10884
rect 3072 10818 3098 10870
rect 3150 10818 3182 10870
rect 3072 10782 3182 10818
rect 3072 10702 3146 10782
rect 3372 10742 3442 10806
rect 3074 10318 3144 10702
rect 3286 10396 3442 10742
rect 3226 10318 3442 10396
rect 3226 10314 3390 10318
rect -9804 10134 -9798 10186
rect -9746 10134 -9740 10186
rect -6772 10160 -6766 10212
rect -6714 10160 -6708 10212
rect -3786 10158 -3780 10210
rect -3728 10158 -3722 10210
rect -778 10156 -772 10208
rect -720 10156 -714 10208
rect 2222 10164 2228 10216
rect 2280 10164 2286 10216
rect 3074 10194 3178 10202
rect 3226 10194 3306 10314
rect 3074 10190 3306 10194
rect 3068 10166 3306 10190
rect 3068 10114 3182 10166
rect 3234 10114 3306 10166
rect 3068 10092 3306 10114
rect 3068 10074 3254 10092
rect 3068 10050 3178 10074
rect 3074 9774 3178 10050
rect 3370 9948 3440 10202
rect 3272 9798 3440 9948
rect -9820 9610 -8742 9754
rect -6808 9608 1916 9748
rect 3250 9738 3440 9798
rect 3250 9606 3298 9738
rect 3370 9714 3440 9738
rect -9650 9326 -8654 9514
rect 3072 9512 3298 9606
rect -6580 9314 -5584 9502
rect -3624 9314 -2628 9502
rect -600 9304 396 9492
rect 3072 9462 3254 9512
rect 3072 9410 3174 9462
rect 3226 9410 3254 9462
rect 3072 9342 3254 9410
rect -11153 9089 -11147 9141
rect -11095 9089 -11089 9141
rect -8154 9124 -8148 9176
rect -8096 9124 -8090 9176
rect -5148 9100 -5142 9152
rect -5090 9100 -5084 9152
rect -2155 9077 -2149 9129
rect -2097 9077 -2091 9129
rect 859 9117 865 9169
rect 917 9117 923 9169
rect 3072 9118 3142 9342
rect 3368 9278 3438 9610
rect 3244 9172 3438 9278
rect 3226 9130 3438 9172
rect 3086 8982 3146 8994
rect 3226 8982 3284 9130
rect 3368 9122 3438 9130
rect 3086 8960 3284 8982
rect 3086 8944 3258 8960
rect 3086 8892 3172 8944
rect 3224 8892 3258 8944
rect 3086 8854 3258 8892
rect 3086 8520 3146 8854
rect 3374 8666 3434 8998
rect 3252 8620 3444 8666
rect 3212 8526 3444 8620
rect 3074 8358 3134 8398
rect 3212 8358 3296 8526
rect 3374 8524 3434 8526
rect 3074 8314 3296 8358
rect 3074 8262 3164 8314
rect 3216 8262 3296 8314
rect 3074 8236 3296 8262
rect 3074 8218 3268 8236
rect 3074 7924 3134 8218
rect 3372 8066 3432 8398
rect 3234 8050 3432 8066
rect 3196 7926 3432 8050
rect 3082 7788 3142 7792
rect 3196 7788 3280 7926
rect 3372 7924 3432 7926
rect 3078 7754 3280 7788
rect 3078 7702 3164 7754
rect 3216 7702 3280 7754
rect 3078 7666 3280 7702
rect 3078 7648 3270 7666
rect -10470 7572 -10464 7624
rect -10412 7572 -10406 7624
rect -7452 7570 -7446 7622
rect -7394 7570 -7388 7622
rect -4454 7556 -4448 7608
rect -4396 7556 -4390 7608
rect -1452 7574 -1446 7626
rect -1394 7574 -1388 7626
rect 1548 7566 1554 7618
rect 1606 7566 1612 7618
rect 3082 7318 3142 7648
rect 3376 7518 3436 7792
rect 3242 7476 3436 7518
rect 3216 7378 3436 7476
rect 3070 7110 3130 7208
rect 3216 7110 3296 7378
rect 3376 7318 3436 7378
rect 3070 7070 3296 7110
rect 3070 7018 3172 7070
rect 3224 7042 3296 7070
rect 3224 7018 3268 7042
rect 3070 6970 3268 7018
rect 3070 6734 3130 6970
rect 3380 6866 3440 7200
rect 3246 6830 3440 6866
rect 3206 6726 3440 6830
rect 3076 6570 3136 6596
rect 3206 6570 3290 6726
rect 3076 6528 3290 6570
rect 3076 6524 3280 6528
rect 3076 6472 3176 6524
rect 3228 6472 3280 6524
rect 3076 6430 3280 6472
rect -9794 6358 -9788 6410
rect -9736 6358 -9730 6410
rect -6792 6348 -6786 6400
rect -6734 6348 -6728 6400
rect -3800 6332 -3794 6384
rect -3742 6332 -3736 6384
rect -778 6330 -772 6382
rect -720 6330 -714 6382
rect 2196 6348 2202 6400
rect 2254 6348 2260 6400
rect 3076 6122 3136 6430
rect 3374 6296 3434 6598
rect 3256 6212 3448 6296
rect 3218 6156 3448 6212
rect 3078 5970 3138 5996
rect 3218 5970 3302 6156
rect 3374 6124 3434 6156
rect -10852 5798 1652 5950
rect 3078 5926 3302 5970
rect 3078 5874 3174 5926
rect 3226 5910 3302 5926
rect 3226 5874 3276 5910
rect 3078 5830 3276 5874
rect -9636 5512 -8640 5700
rect -6656 5504 -5660 5692
rect -3658 5512 -2662 5700
rect -660 5510 336 5698
rect 3078 5522 3138 5830
rect 3370 5680 3430 6000
rect 3244 5648 3436 5680
rect 3208 5540 3436 5648
rect 3208 5398 3292 5540
rect 3370 5526 3430 5540
rect -11146 5296 -11140 5348
rect -11088 5296 -11082 5348
rect -8144 5292 -8138 5344
rect -8086 5292 -8080 5344
rect -5153 5307 -5147 5359
rect -5095 5307 -5089 5359
rect 3078 5358 3292 5398
rect 3078 5306 3174 5358
rect 3226 5346 3292 5358
rect 3226 5306 3270 5346
rect 3078 5258 3270 5306
rect 3080 4918 3140 5258
rect 3370 5090 3430 5408
rect 3248 5016 3440 5090
rect 3222 4950 3440 5016
rect 3080 4766 3140 4806
rect 3222 4766 3306 4950
rect 3370 4934 3430 4950
rect 3072 4718 3306 4766
rect 3072 4666 3178 4718
rect 3230 4714 3306 4718
rect 3230 4666 3264 4714
rect 3072 4626 3264 4666
rect 3080 4332 3140 4626
rect 3374 4468 3434 4802
rect 3240 4446 3434 4468
rect 3202 4328 3434 4446
rect 3074 4202 3134 4210
rect 3202 4202 3286 4328
rect 3074 4150 3286 4202
rect 3074 4098 3176 4150
rect 3228 4144 3286 4150
rect 3228 4098 3266 4144
rect 3074 4062 3266 4098
rect -10460 3762 -10454 3814
rect -10402 3762 -10396 3814
rect -7456 3776 -7450 3828
rect -7398 3776 -7392 3828
rect -4458 3782 -4452 3834
rect -4400 3782 -4394 3834
rect -2162 3734 -2156 3786
rect -2104 3734 -2098 3786
rect -1464 3768 -1458 3820
rect -1406 3768 -1400 3820
rect 837 3794 843 3846
rect 895 3794 901 3846
rect 1558 3790 1564 3842
rect 1616 3790 1622 3842
rect 3074 3736 3134 4062
rect 3378 3924 3438 4208
rect 3234 3840 3438 3924
rect 3202 3784 3438 3840
rect 3074 3522 3134 3604
rect 3202 3522 3284 3784
rect 3378 3734 3438 3784
rect 3074 3492 3284 3522
rect 3074 3440 3178 3492
rect 3230 3476 3284 3492
rect 3230 3440 3270 3476
rect 3074 3382 3270 3440
rect 3074 3130 3134 3382
rect 3370 3272 3430 3604
rect 3236 3216 3430 3272
rect 3236 3204 3296 3216
rect 3210 3158 3296 3204
rect 3352 3158 3430 3216
rect 3210 3132 3430 3158
rect 3210 3006 3272 3132
rect 3370 3130 3430 3132
rect 3072 2954 3272 3006
rect 3072 2866 3264 2954
rect -9762 2578 -9710 2584
rect -6778 2552 -6772 2604
rect -6720 2552 -6714 2604
rect -3778 2562 -3772 2614
rect -3720 2562 -3714 2614
rect -770 2546 -764 2598
rect -712 2546 -706 2598
rect 2178 2576 2378 2582
rect -9762 2520 -9710 2526
rect 3076 2526 3136 2866
rect 3376 2688 3436 3008
rect 3322 2490 3492 2688
rect 2178 2478 2378 2484
rect 2936 2440 3562 2490
rect 2936 2210 2984 2440
rect -10142 1998 1998 2154
rect 2238 2052 2984 2210
rect 3508 2210 3562 2440
rect 3508 2052 3566 2210
rect 2238 2000 3566 2052
<< via1 >>
rect -11152 12894 -11100 12946
rect -8129 12901 -8077 12953
rect -5140 12900 -5088 12952
rect -2129 12903 -2077 12955
rect 3100 12032 3152 12084
rect -10464 11364 -10412 11416
rect -7422 11370 -7370 11422
rect -4434 11364 -4382 11416
rect -1434 11356 -1382 11408
rect 846 11390 898 11442
rect 1552 11374 1604 11426
rect 3098 10818 3150 10870
rect -9798 10134 -9746 10186
rect -6766 10160 -6714 10212
rect -3780 10158 -3728 10210
rect -772 10156 -720 10208
rect 2228 10164 2280 10216
rect 3182 10114 3234 10166
rect 3174 9410 3226 9462
rect -11147 9089 -11095 9141
rect -8148 9124 -8096 9176
rect -5142 9100 -5090 9152
rect -2149 9077 -2097 9129
rect 865 9117 917 9169
rect 3172 8892 3224 8944
rect 3164 8262 3216 8314
rect 3164 7702 3216 7754
rect -10464 7572 -10412 7624
rect -7446 7570 -7394 7622
rect -4448 7556 -4396 7608
rect -1446 7574 -1394 7626
rect 1554 7566 1606 7618
rect 3172 7018 3224 7070
rect 3176 6472 3228 6524
rect -9788 6358 -9736 6410
rect -6786 6348 -6734 6400
rect -3794 6332 -3742 6384
rect -772 6330 -720 6382
rect 2202 6348 2254 6400
rect 3174 5874 3226 5926
rect -11140 5296 -11088 5348
rect -8138 5292 -8086 5344
rect -5147 5307 -5095 5359
rect 3174 5306 3226 5358
rect 3178 4666 3230 4718
rect 3176 4098 3228 4150
rect -10454 3762 -10402 3814
rect -7450 3776 -7398 3828
rect -4452 3782 -4400 3834
rect -2156 3734 -2104 3786
rect -1458 3768 -1406 3820
rect 843 3794 895 3846
rect 1564 3790 1616 3842
rect 3178 3440 3230 3492
rect 3296 3158 3352 3216
rect -9762 2526 -9710 2578
rect -6772 2552 -6720 2604
rect -3772 2562 -3720 2614
rect -764 2546 -712 2598
rect 2178 2484 2378 2576
<< metal2 >>
rect 0 0 100 100
rect 400 0 500 100
rect 1200 0 1300 100
rect 1600 0 1700 100
rect 2000 0 2100 100
rect 2200 0 2300 100
rect 2400 0 2500 100
rect 2600 0 2700 100
rect -5387 13331 2931 13369
rect -5387 13265 -5349 13331
rect -11145 13227 -5349 13265
rect -5274 13261 2853 13302
rect -11145 12952 -11107 13227
rect -5274 13165 -5233 13261
rect -8124 13124 -5233 13165
rect -5129 13183 2765 13213
rect -8124 12959 -8083 13124
rect -8129 12953 -8077 12959
rect -5129 12958 -5099 13183
rect -2124 13097 2677 13138
rect -2124 12961 -2083 13097
rect -11152 12946 -11100 12952
rect -8129 12895 -8077 12901
rect -5140 12952 -5088 12958
rect -5140 12894 -5088 12900
rect -2129 12955 -2077 12961
rect -2129 12897 -2077 12903
rect -11152 12888 -11100 12894
rect 637 11491 1011 11521
rect -13560 11458 -13472 11474
rect -13560 11402 -13542 11458
rect -13486 11402 -13472 11458
rect -7422 11422 -7370 11428
rect -13560 11384 -13472 11402
rect -10464 11416 -10412 11422
rect -16196 11250 -16136 11259
rect -14064 11190 -13614 11218
rect -16196 11181 -16136 11190
rect -13642 10180 -13614 11190
rect -13531 10908 -13496 11384
rect -7422 11364 -7370 11370
rect -4434 11416 -4382 11422
rect -10464 11358 -10412 11364
rect -13404 11248 -13348 11257
rect -13348 11200 -13268 11241
rect -13404 11183 -13348 11192
rect -13531 10873 -13363 10908
rect -13548 10778 -13460 10796
rect -13548 10722 -13532 10778
rect -13476 10722 -13460 10778
rect -13548 10706 -13460 10722
rect -13523 10262 -13484 10706
rect -13398 10346 -13363 10873
rect -13309 10437 -13268 11200
rect -10453 11210 -10423 11358
rect -7411 11231 -7381 11364
rect -4434 11358 -4382 11364
rect -1434 11408 -1382 11414
rect -4423 11231 -4393 11358
rect -1434 11350 -1382 11356
rect -1423 11231 -1393 11350
rect 637 11231 667 11491
rect 846 11442 898 11448
rect 846 11384 898 11390
rect -9225 11210 667 11231
rect -10453 11201 667 11210
rect 858 11206 886 11384
rect 981 11299 1011 11491
rect 1552 11426 1604 11432
rect 1552 11368 1604 11374
rect 1563 11299 1593 11368
rect 981 11269 1593 11299
rect -10453 11180 -9174 11201
rect -13309 10396 -12758 10437
rect -13398 10311 -12839 10346
rect -13523 10223 -12917 10262
rect -13642 10152 -12996 10180
rect -13562 10098 -13474 10118
rect -13562 10042 -13546 10098
rect -13490 10088 -13474 10098
rect -13490 10052 -13070 10088
rect -13490 10042 -13474 10052
rect -13562 10028 -13474 10042
rect -13560 8738 -13472 8760
rect -13560 8682 -13544 8738
rect -13488 8726 -13472 8738
rect -13488 8695 -13157 8726
rect -13488 8682 -13472 8695
rect -13560 8670 -13472 8682
rect -13534 8058 -13442 8072
rect -13534 8002 -13514 8058
rect -13458 8046 -13442 8058
rect -13458 8009 -13237 8046
rect -13458 8002 -13442 8009
rect -13534 7988 -13442 8002
rect -13518 7378 -13426 7386
rect -13518 7322 -13504 7378
rect -13448 7366 -13426 7378
rect -13448 7335 -13325 7366
rect -13448 7322 -13426 7335
rect -13518 7302 -13426 7322
rect -13546 6698 -13458 6712
rect -13546 6642 -13528 6698
rect -13472 6686 -13458 6698
rect -13472 6654 -13398 6686
rect -13472 6642 -13458 6654
rect -13546 6624 -13458 6642
rect -13568 6018 -13480 6034
rect -13568 5962 -13548 6018
rect -13492 5962 -13480 6018
rect -13568 5946 -13480 5962
rect -13674 5338 -13586 5360
rect -13674 5282 -13658 5338
rect -13602 5282 -13586 5338
rect -13674 5272 -13586 5282
rect -14161 2197 -14123 3419
rect -13647 2284 -13612 5272
rect -13537 2366 -13502 5946
rect -13430 5842 -13398 6654
rect -13356 5926 -13325 7335
rect -13274 6001 -13237 8009
rect -13188 6080 -13157 8695
rect -13106 6152 -13070 10052
rect -13024 9758 -12996 10152
rect -12952 9822 -12920 10223
rect -12874 10006 -12839 10311
rect -12799 10077 -12758 10396
rect -6766 10212 -6714 10218
rect -9798 10186 -9746 10192
rect -6766 10154 -6714 10160
rect -3780 10210 -3728 10216
rect -9798 10128 -9746 10134
rect -9793 10077 -9752 10128
rect -12799 10036 -9752 10077
rect -6758 10006 -6723 10154
rect -3780 10152 -3728 10158
rect -772 10208 -720 10214
rect -12874 9971 -6723 10006
rect -12873 9870 -12864 9926
rect -12808 9916 -12799 9926
rect -3772 9916 -3736 10152
rect -772 10150 -720 10156
rect -12808 9880 -3736 9916
rect -12808 9870 -12799 9880
rect -762 9822 -730 10150
rect -111 9897 -81 11201
rect 858 11178 2546 11206
rect 2228 10216 2280 10222
rect 2228 10158 2280 10164
rect -12952 9790 -730 9822
rect -126 9888 -66 9897
rect -126 9819 -66 9828
rect 2240 9758 2268 10158
rect 2518 9794 2546 11178
rect 2636 9902 2677 13097
rect 2735 10145 2765 13183
rect 2812 10822 2853 13261
rect 2893 12069 2931 13331
rect 3080 12084 3174 12108
rect 3080 12069 3100 12084
rect 2893 12032 3100 12069
rect 3152 12032 3174 12084
rect 2893 12031 3174 12032
rect 3080 12008 3174 12031
rect 3082 10870 3176 10884
rect 3082 10822 3098 10870
rect 2812 10818 3098 10822
rect 3150 10818 3176 10870
rect 2812 10784 3176 10818
rect 2812 10781 3149 10784
rect 3164 10166 3258 10186
rect 3164 10145 3182 10166
rect 2735 10115 3182 10145
rect 3164 10114 3182 10115
rect 3234 10114 3258 10166
rect 3164 10086 3258 10114
rect 2636 9861 2985 9902
rect 2518 9766 2878 9794
rect -13024 9730 2268 9758
rect -11141 9642 2806 9681
rect -11141 9147 -11102 9642
rect -8137 9571 2725 9601
rect -8137 9182 -8107 9571
rect -5131 9499 2643 9529
rect -8148 9176 -8096 9182
rect -11147 9141 -11095 9147
rect -5131 9158 -5101 9499
rect -2142 9425 2563 9462
rect -8148 9118 -8096 9124
rect -5142 9152 -5090 9158
rect -2142 9135 -2105 9425
rect 874 9343 2465 9376
rect -126 9184 -66 9186
rect -5142 9094 -5090 9100
rect -2149 9129 -2097 9135
rect -11147 9083 -11095 9089
rect -133 9128 -124 9184
rect -68 9128 -59 9184
rect 874 9175 907 9343
rect 865 9169 917 9175
rect -2149 9071 -2097 9077
rect -10464 7624 -10412 7630
rect -10464 7566 -10412 7572
rect -7446 7622 -7394 7628
rect -1446 7626 -1394 7632
rect -10453 7408 -10423 7566
rect -7446 7564 -7394 7570
rect -4448 7608 -4396 7614
rect -7435 7429 -7405 7564
rect -1446 7568 -1394 7574
rect -4448 7550 -4396 7556
rect -4437 7429 -4407 7550
rect -1435 7429 -1405 7568
rect -126 7464 -66 9128
rect 865 9111 917 9117
rect 1554 7618 1606 7624
rect 1554 7560 1606 7566
rect -220 7429 -66 7464
rect 1565 7429 1595 7560
rect -9293 7408 1595 7429
rect -10453 7399 1595 7408
rect -10453 7378 -9230 7399
rect -220 7344 -66 7399
rect -9788 6410 -9736 6416
rect -9788 6352 -9736 6358
rect -6786 6400 -6734 6406
rect -9780 6152 -9744 6352
rect -3794 6384 -3742 6390
rect -6786 6342 -6734 6348
rect -13106 6116 -9744 6152
rect -6776 6080 -6745 6342
rect -13188 6049 -6745 6080
rect -3797 6332 -3794 6374
rect -3797 6326 -3742 6332
rect -772 6382 -720 6388
rect -3797 6001 -3754 6326
rect -772 6324 -720 6330
rect -13274 5968 -3754 6001
rect -13274 5964 -3760 5968
rect -762 5926 -731 6324
rect -126 6000 -66 7344
rect 2202 6400 2254 6406
rect 2202 6342 2254 6348
rect -126 5931 -66 5940
rect -13356 5895 -731 5926
rect 2212 5842 2244 6342
rect 2432 5919 2465 9343
rect 2526 6491 2563 9425
rect 2613 7059 2643 9499
rect 2695 7743 2725 9571
rect 2767 8306 2806 9642
rect 2850 8932 2878 9766
rect 2944 9459 2985 9861
rect 3158 9462 3252 9490
rect 3158 9459 3174 9462
rect 2944 9418 3174 9459
rect 3158 9410 3174 9418
rect 3226 9410 3252 9462
rect 3158 9390 3252 9410
rect 3156 8944 3250 8966
rect 3156 8932 3172 8944
rect 2850 8904 3172 8932
rect 3156 8892 3172 8904
rect 3224 8892 3250 8944
rect 3156 8866 3250 8892
rect 3148 8314 3242 8344
rect 3148 8306 3164 8314
rect 2767 8267 3164 8306
rect 3148 8262 3164 8267
rect 3216 8262 3242 8314
rect 3148 8244 3242 8262
rect 3144 7754 3238 7782
rect 3144 7743 3164 7754
rect 2695 7713 3164 7743
rect 3144 7702 3164 7713
rect 3216 7702 3238 7754
rect 3144 7682 3238 7702
rect 3154 7070 3248 7094
rect 3154 7059 3172 7070
rect 2613 7029 3172 7059
rect 3154 7018 3172 7029
rect 3224 7018 3248 7070
rect 3154 6994 3248 7018
rect 3154 6524 3248 6556
rect 3154 6491 3176 6524
rect 2526 6472 3176 6491
rect 3228 6472 3248 6524
rect 2526 6456 3248 6472
rect 2526 6454 3184 6456
rect 3158 5926 3252 5952
rect 3158 5919 3174 5926
rect 2432 5886 3174 5919
rect 3158 5874 3174 5886
rect 3226 5919 3252 5926
rect 3226 5886 3256 5919
rect 3226 5874 3252 5886
rect 3158 5852 3252 5874
rect -13430 5810 2244 5842
rect -11131 5735 2675 5769
rect -11131 5354 -11097 5735
rect -8126 5678 2580 5706
rect -11140 5348 -11088 5354
rect -8126 5350 -8098 5678
rect -5141 5576 2472 5615
rect -5141 5365 -5102 5576
rect -126 5440 -66 5442
rect -133 5384 -124 5440
rect -68 5384 -59 5440
rect -5147 5359 -5095 5365
rect -11140 5290 -11088 5296
rect -8138 5344 -8086 5350
rect -5147 5301 -5095 5307
rect -8138 5286 -8086 5292
rect -13454 4658 -13366 4680
rect -13454 4602 -13442 4658
rect -13386 4602 -13366 4658
rect -13454 4592 -13366 4602
rect -13434 2473 -13393 4592
rect -13318 3978 -13262 3987
rect -13318 3913 -13262 3922
rect -2311 3951 -2001 3981
rect -13309 2571 -13271 3913
rect -4452 3834 -4400 3840
rect -7450 3828 -7398 3834
rect -10454 3814 -10402 3820
rect -4452 3776 -4400 3782
rect -7450 3770 -7398 3776
rect -10454 3756 -10402 3762
rect -10443 3626 -10413 3756
rect -7439 3626 -7409 3770
rect -4441 3626 -4411 3776
rect -2311 3626 -2281 3951
rect -2156 3786 -2104 3792
rect -2156 3728 -2104 3734
rect -10443 3596 -2281 3626
rect -2150 3624 -2110 3728
rect -2031 3713 -2001 3951
rect -1458 3820 -1406 3826
rect -1406 3768 -1390 3806
rect -1458 3762 -1390 3768
rect -1447 3740 -1390 3762
rect -1447 3735 -156 3740
rect -126 3735 -66 5384
rect 2433 4142 2472 5576
rect 2552 4708 2580 5678
rect 2641 5343 2675 5735
rect 3140 5358 3252 5372
rect 3140 5343 3174 5358
rect 2641 5309 3174 5343
rect 3140 5306 3174 5309
rect 3226 5306 3252 5358
rect 3140 5282 3252 5306
rect 3150 4718 3262 4734
rect 3150 4708 3178 4718
rect 2552 4680 3178 4708
rect 3150 4666 3178 4680
rect 3230 4666 3262 4718
rect 3150 4644 3262 4666
rect 3140 4150 3252 4168
rect 3140 4142 3176 4150
rect 2433 4103 3176 4142
rect 3140 4098 3176 4103
rect 3228 4098 3252 4150
rect 3140 4078 3252 4098
rect 539 4034 1041 4041
rect 539 3999 1046 4034
rect 539 3735 581 3999
rect -1447 3713 581 3735
rect -2031 3693 581 3713
rect 774 3902 982 3942
rect -2031 3688 -156 3693
rect -2031 3683 -1417 3688
rect 774 3624 814 3902
rect 843 3846 895 3852
rect 843 3788 895 3794
rect -2150 3584 814 3624
rect 848 3582 889 3788
rect 942 3660 982 3902
rect 1018 3734 1046 3999
rect 1564 3842 1616 3848
rect 1564 3784 1616 3790
rect 1576 3734 1604 3784
rect 1018 3706 1604 3734
rect 942 3620 2536 3660
rect 848 3541 2439 3582
rect 2398 3207 2439 3541
rect 2496 3482 2536 3620
rect 3138 3492 3250 3508
rect 3138 3482 3178 3492
rect 2496 3442 3178 3482
rect 3138 3440 3178 3442
rect 3230 3440 3250 3492
rect 3138 3418 3250 3440
rect 3274 3216 3368 3226
rect 3274 3207 3296 3216
rect 2398 3166 3296 3207
rect 3274 3158 3296 3166
rect 3352 3158 3368 3216
rect 3274 3142 3368 3158
rect -3772 2614 -3720 2620
rect -6772 2604 -6720 2610
rect -9768 2571 -9762 2578
rect -13309 2533 -9762 2571
rect -9768 2526 -9762 2533
rect -9710 2526 -9704 2578
rect -3772 2556 -3720 2562
rect -764 2598 -712 2604
rect -6772 2546 -6720 2552
rect -6767 2473 -6726 2546
rect -13434 2432 -6726 2473
rect -3764 2366 -3729 2556
rect -764 2540 -712 2546
rect -13537 2331 -3729 2366
rect -756 2284 -721 2540
rect 2172 2484 2178 2576
rect 2378 2484 2384 2576
rect -13647 2249 -721 2284
rect 2259 2197 2297 2484
rect -14161 2159 2297 2197
<< via2 >>
rect -13542 11402 -13486 11458
rect -16196 11190 -16136 11250
rect -13404 11192 -13348 11248
rect -13532 10722 -13476 10778
rect -13546 10042 -13490 10098
rect -13544 8682 -13488 8738
rect -13514 8002 -13458 8058
rect -13504 7322 -13448 7378
rect -13528 6642 -13472 6698
rect -13548 5962 -13492 6018
rect -13658 5282 -13602 5338
rect -12864 9870 -12808 9926
rect -126 9828 -66 9888
rect -124 9128 -68 9184
rect -126 5940 -66 6000
rect -124 5384 -68 5440
rect -13442 4602 -13386 4658
rect -13318 3922 -13262 3978
<< metal3 >>
rect 200 0 300 100
rect 600 0 700 100
rect 1400 0 1500 100
rect 1800 0 1900 100
rect 2800 0 2900 100
rect -13560 11458 -13472 11474
rect -13560 11402 -13542 11458
rect -13486 11402 -13472 11458
rect -13560 11384 -13472 11402
rect -16201 11250 -16131 11255
rect -13409 11250 -13343 11253
rect -16201 11190 -16196 11250
rect -16136 11248 -13343 11250
rect -16136 11192 -13404 11248
rect -13348 11192 -13343 11248
rect -16136 11190 -13343 11192
rect -16201 11185 -16131 11190
rect -13409 11187 -13343 11190
rect -13548 10778 -13460 10796
rect -13548 10722 -13532 10778
rect -13476 10722 -13460 10778
rect -13548 10706 -13460 10722
rect -13562 10098 -13474 10118
rect -13562 10042 -13546 10098
rect -13490 10042 -13474 10098
rect -13562 10028 -13474 10042
rect -12869 9926 -12803 9931
rect -12869 9870 -12864 9926
rect -12808 9870 -12803 9926
rect -12869 9865 -12803 9870
rect -131 9888 -61 9893
rect -12866 9420 -12806 9865
rect -131 9828 -126 9888
rect -66 9828 -61 9888
rect -131 9823 -61 9828
rect -13534 9360 -12806 9420
rect -126 9189 -66 9823
rect -129 9184 -63 9189
rect -129 9128 -124 9184
rect -68 9128 -63 9184
rect -129 9123 -63 9128
rect -13560 8738 -13472 8760
rect -13560 8682 -13544 8738
rect -13488 8682 -13472 8738
rect -13560 8670 -13472 8682
rect -13470 8078 -13364 8090
rect -13534 8058 -13364 8078
rect -13534 8002 -13514 8058
rect -13458 8002 -13364 8058
rect -13534 7988 -13364 8002
rect -13470 7978 -13364 7988
rect -13450 7386 -13374 7400
rect -13518 7378 -13374 7386
rect -13518 7322 -13504 7378
rect -13448 7322 -13374 7378
rect -13518 7302 -13374 7322
rect -13450 7292 -13374 7302
rect -13478 6712 -13382 6722
rect -13546 6698 -13382 6712
rect -13546 6642 -13528 6698
rect -13472 6642 -13382 6698
rect -13546 6624 -13382 6642
rect -13478 6610 -13382 6624
rect -13568 6018 -13480 6034
rect -13568 5962 -13548 6018
rect -13492 5962 -13480 6018
rect -13568 5946 -13480 5962
rect -131 6000 -61 6005
rect -131 5940 -126 6000
rect -66 5940 -61 6000
rect -131 5935 -61 5940
rect -126 5445 -66 5935
rect -129 5440 -63 5445
rect -129 5384 -124 5440
rect -68 5384 -63 5440
rect -129 5379 -63 5384
rect -13674 5338 -13586 5360
rect -13674 5282 -13658 5338
rect -13602 5282 -13586 5338
rect -13674 5272 -13586 5282
rect -13454 4658 -13366 4680
rect -13454 4602 -13442 4658
rect -13386 4602 -13366 4658
rect -13454 4592 -13366 4602
rect -13316 3983 -12950 3984
rect -13323 3978 -12950 3983
rect -13323 3922 -13318 3978
rect -13262 3922 -12950 3978
rect -13323 3917 -12950 3922
rect -13316 3916 -12950 3917
<< metal4 >>
rect 0 0 100 100 0
rect 200 0 300 100 0
rect 400 0 500 100 0
rect 600 0 700 100 0


use bit4_encoder  bit4_encoder_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730718415
transform 1 0 -22008 0 1 1842
box 0 0 9409 11553
use compr  compr_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730635755
transform 1 0 -1234 0 1 2394
box 1230 -398 4034 3312
use compr  compr_1
timestamp 1730635755
transform 1 0 -4232 0 1 2394
box 1230 -398 4034 3312
use compr  compr_2
timestamp 1730635755
transform 1 0 -7238 0 1 2394
box 1230 -398 4034 3312
use compr  compr_3
timestamp 1730635755
transform 1 0 -10234 0 1 2394
box 1230 -398 4034 3312
use compr  compr_4
timestamp 1730635755
transform 1 0 -13232 0 1 2394
box 1230 -398 4034 3312
use compr  compr_5
timestamp 1730635755
transform 1 0 -1230 0 1 6192
box 1230 -398 4034 3312
use compr  compr_6
timestamp 1730635755
transform 1 0 -4226 0 1 6192
box 1230 -398 4034 3312
use compr  compr_7
timestamp 1730635755
transform 1 0 -7230 0 1 6192
box 1230 -398 4034 3312
use compr  compr_8
timestamp 1730635755
transform 1 0 -10234 0 1 6202
box 1230 -398 4034 3312
use compr  compr_9
timestamp 1730635755
transform 1 0 -13238 0 1 6202
box 1230 -398 4034 3312
use compr  compr_10
timestamp 1730635755
transform 1 0 -1230 0 1 10002
box 1230 -398 4034 3312
use compr  compr_11
timestamp 1730635755
transform 1 0 -4226 0 1 9992
box 1230 -398 4034 3312
use compr  compr_12
timestamp 1730635755
transform 1 0 -7230 0 1 9992
box 1230 -398 4034 3312
use compr  compr_13
timestamp 1730635755
transform 1 0 -10234 0 1 10002
box 1230 -398 4034 3312
use compr  compr_14
timestamp 1730635755
transform 1 0 -13246 0 1 9992
box 1230 -398 4034 3312
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR1
timestamp 1730493024
transform 1 0 3107 0 1 11458
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730493024
transform 1 0 3403 0 1 6666
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR3
timestamp 1730493024
transform 1 0 3403 0 1 10260
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR4
timestamp 1730493024
transform 1 0 3107 0 1 12656
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR5
timestamp 1730493024
transform 1 0 3403 0 1 7864
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730493024
transform 1 0 3107 0 1 3072
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR7
timestamp 1730493024
transform 1 0 3403 0 1 9062
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730493024
transform 1 0 3107 0 1 5468
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR9
timestamp 1730493024
transform 1 0 3107 0 1 10260
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730493024
transform 1 0 3107 0 1 6666
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR11
timestamp 1730493024
transform 1 0 3107 0 1 9062
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730493024
transform 1 0 3107 0 1 7864
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR13
timestamp 1730493024
transform 1 0 3403 0 1 3072
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730493024
transform 1 0 3403 0 1 4270
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR15
timestamp 1730493024
transform 1 0 3403 0 1 5468
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730493024
transform 1 0 3107 0 1 4270
box -201 -652 201 652
<< labels >>
flabel metal2 s 0 0 100 100 0 FreeSans 480 90 0 0 bus00
port 0 nsew
flabel metal3 s 200 0 300 100 0 FreeSans 480 90 0 0 bus01
port 1 nsew
flabel metal2 s 400 0 500 100 0 FreeSans 480 90 0 0 bus02
port 2 nsew
flabel metal3 s 600 0 700 100 0 FreeSans 480 90 0 0 bus03
port 3 nsew
flabel metal2 s 1200 0 1300 100 0 FreeSans 480 90 0 0 bus10
port 4 nsew
flabel metal3 s 1400 0 1500 100 0 FreeSans 480 90 0 0 bus11
port 5 nsew
flabel metal2 s 1600 0 1700 100 0 FreeSans 480 90 0 0 bus12
port 6 nsew
flabel metal3 s 1800 0 1900 100 0 FreeSans 480 90 0 0 bus13
port 7 nsew
flabel metal2 s 2000 0 2100 100 0 FreeSans 480 90 0 0 bus20
port 8 nsew
flabel metal2 s 2200 0 2300 100 0 FreeSans 480 90 0 0 bus21
port 9 nsew
flabel metal2 s 2400 0 2500 100 0 FreeSans 480 90 0 0 bus22
port 10 nsew
flabel metal2 s 2600 0 2700 100 0 FreeSans 480 90 0 0 bus23
port 11 nsew
flabel metal3 s 2800 0 2900 100 0 FreeSans 480 90 0 0 clk
port 12 nsew
flabel metal1 800 0 900 100 1 FreeSans 400 0 0 0 VDPWR
port 13 nsew power bidirectional
flabel metal1 1000 0 1100 100 1 FreeSans 400 0 0 0 VGND
port 14 nsew ground bidirectional
<< end >>
