* NGSPICE file created from variable_delay_dummy_parax.ext - technology: sky130A

.subckt variable_delay_dummy_parax in out VSS VDD
X0 VDD.t36 VDD.t34 a_5444_772# VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1 VDD.t33 VDD.t31 a_2496_772# VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X2 VDD.t30 VDD.t28 a_5444_772# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X3 VSS.t33 variable_delay_unit_1.tristate_inverter_1.en.t2 a_5444_352# VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X4 variable_delay_unit_1.out variable_delay_unit_1.forward.t2 a_4562_772# VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X5 VSS.t35 variable_delay_unit_0.tristate_inverter_1.en.t2 a_2496_352# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X6 VSS.t31 variable_delay_unit_1.tristate_inverter_1.en.t3 a_5444_352# VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X7 variable_delay_unit_0.tristate_inverter_1.en.t1 VDD.t25 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X8 VDD.t43 variable_delay_unit_1.tristate_inverter_1.en.t4 a_4562_772# VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X9 out.t3 variable_delay_unit_1.in.t2 a_1614_772# VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X10 VSS.t24 VDD.t44 a_4562_352# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 variable_delay_unit_1.out variable_delay_unit_1.forward.t3 a_4562_352# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X12 variable_delay_unit_0.tristate_inverter_1.en.t0 VDD.t45 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X13 out.t2 variable_delay_unit_1.in.t3 a_1614_352# VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X14 a_2496_772# variable_delay_unit_1.out out.t0 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X15 a_2496_352# variable_delay_unit_1.out out.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X16 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t3 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X17 a_5444_772# VDD.t22 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X18 a_1614_352# VDD.t46 VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X19 variable_delay_unit_1.tristate_inverter_1.en.t1 VDD.t19 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X20 a_5444_772# VSS.t37 variable_delay_unit_1.out VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X21 variable_delay_unit_1.tristate_inverter_1.en.t0 VDD.t47 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X22 a_5444_352# variable_delay_unit_1.tristate_inverter_1.en.t5 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X23 a_2496_772# VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X24 a_2496_352# variable_delay_unit_0.tristate_inverter_1.en.t4 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X25 a_5444_352# VSS.t2 variable_delay_unit_1.out VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X26 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t5 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X27 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t6 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X28 a_1614_352# VDD.t48 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X29 a_4562_352# VDD.t49 VSS.t14 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X30 variable_delay_unit_1.in.t0 in.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X31 variable_delay_unit_1.in.t1 in.t1 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X32 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t7 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X33 a_4562_352# VDD.t50 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X34 VDD.t15 VDD.t13 a_2496_772# VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X35 variable_delay_unit_1.forward.t1 variable_delay_unit_1.in.t4 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X36 VSS.t7 variable_delay_unit_0.tristate_inverter_1.en.t6 a_2496_352# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X37 variable_delay_unit_1.forward.t0 variable_delay_unit_1.in.t5 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X38 VDD.t7 variable_delay_unit_0.tristate_inverter_1.en.t7 a_1614_772# VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X39 VSS.t10 VDD.t51 a_1614_352# VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
R0 VDD.n106 VDD.n64 1689.71
R1 VDD.n69 VDD.n64 1689.71
R2 VDD.n62 VDD.n61 1689.71
R3 VDD.n109 VDD.n61 1689.71
R4 VDD.n30 VDD.n13 1689.71
R5 VDD.n30 VDD.n14 1689.71
R6 VDD.n20 VDD.n15 1689.71
R7 VDD.n26 VDD.n15 1689.71
R8 VDD.n44 VDD.n3 1307.92
R9 VDD.n40 VDD.n4 1307.92
R10 VDD.n89 VDD.n77 1307.92
R11 VDD.n74 VDD.n73 1307.92
R12 VDD.n79 VDD.t31 628.097
R13 VDD.n50 VDD.t34 628.097
R14 VDD.n80 VDD.t13 622.766
R15 VDD.n51 VDD.t28 622.766
R16 VDD.n83 VDD.t25 543.053
R17 VDD.n54 VDD.t19 543.053
R18 VDD.n79 VDD.t16 523.774
R19 VDD.n50 VDD.t22 523.774
R20 VDD.n108 VDD.n107 332.803
R21 VDD.n28 VDD.n27 332.803
R22 VDD.n78 VDD.t46 304.647
R23 VDD.n78 VDD.t48 304.647
R24 VDD.n49 VDD.t49 304.647
R25 VDD.n49 VDD.t50 304.647
R26 VDD.n83 VDD.t45 221.72
R27 VDD.n54 VDD.t47 221.72
R28 VDD.n84 VDD.n83 219.549
R29 VDD.n55 VDD.n54 219.531
R30 VDD.n78 VDD.t51 202.44
R31 VDD.n49 VDD.t44 202.44
R32 VDD.n105 VDD.n65 180.236
R33 VDD.n70 VDD.n65 180.236
R34 VDD.n111 VDD.n110 180.236
R35 VDD.n111 VDD.n57 180.236
R36 VDD.n31 VDD.n12 180.236
R37 VDD.n31 VDD.n8 180.236
R38 VDD.n25 VDD.n16 180.236
R39 VDD.n21 VDD.n16 180.236
R40 VDD.n43 VDD.n0 175.123
R41 VDD.n7 VDD.n6 175.123
R42 VDD.n92 VDD.n91 175.123
R43 VDD.n87 VDD.n71 175.123
R44 VDD VDD.n78 168.969
R45 VDD VDD.n49 168.969
R46 VDD VDD.n80 166.147
R47 VDD VDD.n51 166.147
R48 VDD.t32 VDD.n62 163.724
R49 VDD.n69 VDD.t1 163.724
R50 VDD.n20 VDD.t35 163.724
R51 VDD.t9 VDD.n14 163.724
R52 VDD.n41 VDD.t37 160.923
R53 VDD.t20 VDD.n42 160.923
R54 VDD.n88 VDD.t4 160.923
R55 VDD.t26 VDD.n90 160.923
R56 VDD.n108 VDD.t8 145.224
R57 VDD.n107 VDD.t3 145.224
R58 VDD.n27 VDD.t0 145.224
R59 VDD.t39 VDD.n28 145.224
R60 VDD.n45 VDD.n2 139.512
R61 VDD.n45 VDD.n0 139.512
R62 VDD.n39 VDD.n5 139.512
R63 VDD.n7 VDD.n5 139.512
R64 VDD.n93 VDD.n75 139.512
R65 VDD.n93 VDD.n92 139.512
R66 VDD.n98 VDD.n97 139.512
R67 VDD.n98 VDD.n71 139.512
R68 VDD.n42 VDD.n41 119.861
R69 VDD.n90 VDD.n88 119.861
R70 VDD.t17 VDD.t32 88.7478
R71 VDD.t8 VDD.t14 88.7478
R72 VDD.t11 VDD.t3 88.7478
R73 VDD.t1 VDD.t6 88.7478
R74 VDD.t35 VDD.t23 88.7478
R75 VDD.t29 VDD.t0 88.7478
R76 VDD.t40 VDD.t39 88.7478
R77 VDD.t42 VDD.t9 88.7478
R78 VDD.n47 VDD.t21 84.7934
R79 VDD.n37 VDD.t38 84.7934
R80 VDD.n76 VDD.t27 84.7934
R81 VDD.n72 VDD.t5 84.7934
R82 VDD.n67 VDD.n66 84.7744
R83 VDD.n59 VDD.n58 84.7744
R84 VDD.n10 VDD.n9 84.7744
R85 VDD.n18 VDD.n17 84.7744
R86 VDD.n67 VDD.t2 83.8097
R87 VDD.n59 VDD.t33 83.8097
R88 VDD.n10 VDD.t10 83.8097
R89 VDD.n18 VDD.t36 83.8097
R90 VDD.n45 VDD.n44 46.2505
R91 VDD.n5 VDD.n4 46.2505
R92 VDD.n93 VDD.n77 46.2505
R93 VDD.n98 VDD.n73 46.2505
R94 VDD.n63 VDD.t17 44.3742
R95 VDD.t14 VDD.n63 44.3742
R96 VDD.n68 VDD.t11 44.3742
R97 VDD.t6 VDD.n68 44.3742
R98 VDD.t23 VDD.n19 44.3742
R99 VDD.n19 VDD.t29 44.3742
R100 VDD.n29 VDD.t40 44.3742
R101 VDD.n29 VDD.t42 44.3742
R102 VDD.n44 VDD.n43 39.3924
R103 VDD.n6 VDD.n4 39.3924
R104 VDD.n91 VDD.n77 39.3924
R105 VDD.n87 VDD.n73 39.3924
R106 VDD.n65 VDD.n64 23.1255
R107 VDD.n68 VDD.n64 23.1255
R108 VDD.n111 VDD.n61 23.1255
R109 VDD.n63 VDD.n61 23.1255
R110 VDD.n31 VDD.n30 23.1255
R111 VDD.n30 VDD.n29 23.1255
R112 VDD.n16 VDD.n15 23.1255
R113 VDD.n19 VDD.n15 23.1255
R114 VDD.n3 VDD.n2 20.5561
R115 VDD.n42 VDD.n3 20.5561
R116 VDD.n40 VDD.n39 20.5561
R117 VDD.n41 VDD.n40 20.5561
R118 VDD.n89 VDD.n75 20.5561
R119 VDD.n90 VDD.n89 20.5561
R120 VDD.n97 VDD.n74 20.5561
R121 VDD.n88 VDD.n74 20.5561
R122 VDD.n70 VDD.n69 18.5005
R123 VDD.n106 VDD.n105 18.5005
R124 VDD.n107 VDD.n106 18.5005
R125 VDD.n110 VDD.n109 18.5005
R126 VDD.n109 VDD.n108 18.5005
R127 VDD.n62 VDD.n57 18.5005
R128 VDD.n14 VDD.n8 18.5005
R129 VDD.n13 VDD.n12 18.5005
R130 VDD.n28 VDD.n13 18.5005
R131 VDD.n26 VDD.n25 18.5005
R132 VDD.n27 VDD.n26 18.5005
R133 VDD.n21 VDD.n20 18.5005
R134 VDD.n66 VDD.t12 9.52217
R135 VDD.n66 VDD.t7 9.52217
R136 VDD.n58 VDD.t18 9.52217
R137 VDD.n58 VDD.t15 9.52217
R138 VDD.n9 VDD.t41 9.52217
R139 VDD.n9 VDD.t43 9.52217
R140 VDD.n17 VDD.t24 9.52217
R141 VDD.n17 VDD.t30 9.52217
R142 VDD.n6 VDD.t37 5.4667
R143 VDD.n43 VDD.t20 5.4667
R144 VDD.t4 VDD.n87 5.4667
R145 VDD.n91 VDD.t26 5.4667
R146 VDD.n82 VDD.n81 3.26479
R147 VDD.n53 VDD.n52 3.26479
R148 VDD.n36 VDD.n5 2.3255
R149 VDD.n46 VDD.n45 2.3255
R150 VDD.n99 VDD.n98 2.3255
R151 VDD.n94 VDD.n93 2.3255
R152 VDD.n56 VDD.n55 2.2505
R153 VDD.n85 VDD.n84 2.2505
R154 VDD.n39 VDD.n38 2.04321
R155 VDD.n48 VDD.n0 2.04321
R156 VDD.n2 VDD.n1 2.04321
R157 VDD.n35 VDD.n7 2.04321
R158 VDD.n97 VDD.n96 2.04321
R159 VDD.n92 VDD.n86 2.04321
R160 VDD.n95 VDD.n75 2.04321
R161 VDD.n100 VDD.n71 2.04321
R162 VDD VDD.n21 1.97234
R163 VDD.n110 VDD.n60 1.96583
R164 VDD.n101 VDD.n70 1.96583
R165 VDD.n105 VDD.n104 1.96583
R166 VDD.n114 VDD.n57 1.96583
R167 VDD.n25 VDD.n24 1.96583
R168 VDD.n34 VDD.n8 1.96583
R169 VDD.n12 VDD.n11 1.96583
R170 VDD.n81 VDD 1.40175
R171 VDD.n52 VDD 1.40175
R172 VDD.n23 VDD.n16 1.32907
R173 VDD.n32 VDD.n31 1.32907
R174 VDD.n112 VDD.n111 1.32907
R175 VDD.n103 VDD.n65 1.32907
R176 VDD.n102 VDD.n67 1.21789
R177 VDD.n113 VDD.n59 1.21789
R178 VDD.n33 VDD.n10 1.21789
R179 VDD.n22 VDD.n18 1.21789
R180 VDD.n80 VDD.n79 1.09595
R181 VDD.n51 VDD.n50 1.09595
R182 VDD.n55 VDD.n53 0.732643
R183 VDD.n84 VDD.n82 0.714786
R184 VDD.n81 VDD 0.443357
R185 VDD.n52 VDD 0.443357
R186 VDD.n35 VDD 0.432792
R187 VDD VDD.n100 0.432792
R188 VDD.n24 VDD.n11 0.430188
R189 VDD.n104 VDD.n60 0.430188
R190 VDD VDD.n56 0.385917
R191 VDD.n24 VDD.n23 0.359875
R192 VDD.n32 VDD.n11 0.359875
R193 VDD.n112 VDD.n60 0.359875
R194 VDD.n104 VDD.n103 0.359875
R195 VDD.n85 VDD 0.297375
R196 VDD.n23 VDD.n22 0.229667
R197 VDD.n33 VDD.n32 0.229667
R198 VDD.n113 VDD.n112 0.229667
R199 VDD.n103 VDD.n102 0.229667
R200 VDD.n86 VDD.n85 0.195812
R201 VDD.n36 VDD.n35 0.189302
R202 VDD.n46 VDD.n1 0.189302
R203 VDD.n100 VDD.n99 0.189302
R204 VDD.n95 VDD.n94 0.189302
R205 VDD.n56 VDD.n48 0.182792
R206 VDD.n38 VDD.n1 0.141125
R207 VDD.n96 VDD.n95 0.141125
R208 VDD.n38 VDD.n37 0.13201
R209 VDD.n48 VDD.n47 0.13201
R210 VDD.n96 VDD.n72 0.13201
R211 VDD.n86 VDD.n76 0.13201
R212 VDD.n34 VDD.n33 0.130708
R213 VDD.n102 VDD.n101 0.130708
R214 VDD.n22 VDD 0.124198
R215 VDD VDD.n113 0.124198
R216 VDD VDD.n34 0.0695104
R217 VDD VDD.n114 0.0695104
R218 VDD.n101 VDD 0.0695104
R219 VDD.n82 VDD 0.063
R220 VDD.n53 VDD 0.063
R221 VDD.n37 VDD.n36 0.0577917
R222 VDD.n47 VDD.n46 0.0577917
R223 VDD.n99 VDD.n72 0.0577917
R224 VDD.n94 VDD.n76 0.0577917
R225 VDD.n114 VDD 0.00701042
R226 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t6 628.097
R227 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.t7 622.766
R228 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t4 523.774
R229 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t3 304.647
R230 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t2 304.647
R231 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t5 202.44
R232 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n0 168.969
R233 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n4 166.147
R234 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t1 84.7557
R235 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t0 84.1197
R236 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R237 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en 5.58443
R238 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n2 4.59003
R239 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.n3 1.09595
R240 VSS.n77 VSS.n76 50016.6
R241 VSS.n85 VSS.n78 23663.9
R242 VSS.n86 VSS.n85 22860.5
R243 VSS.n77 VSS.n21 14239.4
R244 VSS.n85 VSS.n84 14239.4
R245 VSS.n78 VSS.n77 10823.2
R246 VSS.n78 VSS.n20 10102.8
R247 VSS.n64 VSS.n63 2045.07
R248 VSS.n109 VSS.n108 2045.07
R249 VSS.n110 VSS.n5 1626.7
R250 VSS.n18 VSS.n5 1626.7
R251 VSS.n67 VSS.n61 1626.7
R252 VSS.n67 VSS.n60 1626.7
R253 VSS.n29 VSS.n22 1626.7
R254 VSS.n75 VSS.n22 1626.7
R255 VSS.n80 VSS.n6 1626.7
R256 VSS.n107 VSS.n6 1626.7
R257 VSS.n44 VSS.n20 1460.78
R258 VSS.n20 VSS.n19 1437.75
R259 VSS.n39 VSS.n21 1138.52
R260 VSS.n84 VSS.n83 1138.52
R261 VSS.n65 VSS.n21 1115.49
R262 VSS.n84 VSS.n81 1115.49
R263 VSS.n45 VSS.n40 1058.19
R264 VSS.n51 VSS.n40 1058.19
R265 VSS.n54 VSS.n38 1058.19
R266 VSS.n54 VSS.n37 1058.19
R267 VSS.n87 VSS.n15 1058.19
R268 VSS.n94 VSS.n15 1058.19
R269 VSS.n97 VSS.n13 1058.19
R270 VSS.n82 VSS.n13 1058.19
R271 VSS.t25 VSS.n39 943.788
R272 VSS.t25 VSS.n53 943.788
R273 VSS.n52 VSS.t17 943.788
R274 VSS.n44 VSS.t17 943.788
R275 VSS.n83 VSS.t4 943.788
R276 VSS.n96 VSS.t4 943.788
R277 VSS.n95 VSS.t19 943.788
R278 VSS.n86 VSS.t19 943.788
R279 VSS.n76 VSS.t32 892.394
R280 VSS.n63 VSS.t3 892.394
R281 VSS.t27 VSS.n64 892.394
R282 VSS.t13 VSS.n65 892.394
R283 VSS.n19 VSS.t34 892.394
R284 VSS.n109 VSS.t8 892.394
R285 VSS.n108 VSS.t36 892.394
R286 VSS.n81 VSS.t21 892.394
R287 VSS.n53 VSS.n52 702.96
R288 VSS.n96 VSS.n95 702.96
R289 VSS.n23 VSS.t37 607.409
R290 VSS.t28 VSS.t32 545.352
R291 VSS.t3 VSS.t30 545.352
R292 VSS.t11 VSS.t27 545.352
R293 VSS.t23 VSS.t13 545.352
R294 VSS.t34 VSS.t0 545.352
R295 VSS.t6 VSS.t8 545.352
R296 VSS.t15 VSS.t36 545.352
R297 VSS.t21 VSS.t9 545.352
R298 VSS.n23 VSS.t2 321.423
R299 VSS.n62 VSS.t28 272.676
R300 VSS.t30 VSS.n62 272.676
R301 VSS.n66 VSS.t11 272.676
R302 VSS.n66 VSS.t23 272.676
R303 VSS.t0 VSS.n17 272.676
R304 VSS.n17 VSS.t6 272.676
R305 VSS.n79 VSS.t15 272.676
R306 VSS.t9 VSS.n79 272.676
R307 VSS.n37 VSS.n34 195
R308 VSS.n39 VSS.n37 195
R309 VSS.n38 VSS.n36 195
R310 VSS.n53 VSS.n38 195
R311 VSS.n51 VSS.n50 195
R312 VSS.n52 VSS.n51 195
R313 VSS.n48 VSS.n45 195
R314 VSS.n45 VSS.n44 195
R315 VSS.n82 VSS.n11 195
R316 VSS.n83 VSS.n82 195
R317 VSS.n98 VSS.n97 195
R318 VSS.n97 VSS.n96 195
R319 VSS.n94 VSS.n93 195
R320 VSS.n95 VSS.n94 195
R321 VSS.n88 VSS.n87 195
R322 VSS.n87 VSS.n86 195
R323 VSS VSS.n23 161.595
R324 VSS.n55 VSS.n54 146.25
R325 VSS.n54 VSS.t25 146.25
R326 VSS.n49 VSS.n40 146.25
R327 VSS.n40 VSS.t17 146.25
R328 VSS.n75 VSS.n74 146.25
R329 VSS.n76 VSS.n75 146.25
R330 VSS.n72 VSS.n29 146.25
R331 VSS.n63 VSS.n29 146.25
R332 VSS.n60 VSS.n30 146.25
R333 VSS.n64 VSS.n60 146.25
R334 VSS.n61 VSS.n59 146.25
R335 VSS.n65 VSS.n61 146.25
R336 VSS.n99 VSS.n13 146.25
R337 VSS.t4 VSS.n13 146.25
R338 VSS.n92 VSS.n15 146.25
R339 VSS.n15 VSS.t19 146.25
R340 VSS.n18 VSS.n4 146.25
R341 VSS.n19 VSS.n18 146.25
R342 VSS.n111 VSS.n110 146.25
R343 VSS.n110 VSS.n109 146.25
R344 VSS.n107 VSS.n106 146.25
R345 VSS.n108 VSS.n107 146.25
R346 VSS.n80 VSS.n10 146.25
R347 VSS.n81 VSS.n80 146.25
R348 VSS.n112 VSS.n111 105.695
R349 VSS.n112 VSS.n4 105.695
R350 VSS.n74 VSS.n73 105.695
R351 VSS.n73 VSS.n72 105.695
R352 VSS.n68 VSS.n30 105.695
R353 VSS.n68 VSS.n59 105.695
R354 VSS.n106 VSS.n7 105.695
R355 VSS.n10 VSS.n7 105.695
R356 VSS.n12 VSS.t5 84.1574
R357 VSS.n90 VSS.t20 84.1574
R358 VSS.n35 VSS.t26 84.1574
R359 VSS.n46 VSS.t18 84.1574
R360 VSS.n2 VSS.t35 83.7172
R361 VSS.n9 VSS.t22 83.7172
R362 VSS.n26 VSS.t33 83.7172
R363 VSS.n32 VSS.t14 83.7172
R364 VSS.n2 VSS.n1 75.905
R365 VSS.n9 VSS.n8 75.905
R366 VSS.n26 VSS.n25 75.905
R367 VSS.n32 VSS.n31 75.905
R368 VSS.n73 VSS.n22 73.1255
R369 VSS.n62 VSS.n22 73.1255
R370 VSS.n68 VSS.n67 73.1255
R371 VSS.n67 VSS.n66 73.1255
R372 VSS.n112 VSS.n5 73.1255
R373 VSS.n17 VSS.n5 73.1255
R374 VSS.n7 VSS.n6 73.1255
R375 VSS.n79 VSS.n6 73.1255
R376 VSS.n50 VSS.n49 68.7561
R377 VSS.n49 VSS.n48 68.7561
R378 VSS.n55 VSS.n36 68.7561
R379 VSS.n55 VSS.n34 68.7561
R380 VSS.n92 VSS.n88 68.7561
R381 VSS.n93 VSS.n92 68.7561
R382 VSS.n99 VSS.n98 68.7561
R383 VSS.n99 VSS.n11 68.7561
R384 VSS.n1 VSS.t1 17.4005
R385 VSS.n1 VSS.t7 17.4005
R386 VSS.n8 VSS.t16 17.4005
R387 VSS.n8 VSS.t10 17.4005
R388 VSS.n25 VSS.t29 17.4005
R389 VSS.n25 VSS.t31 17.4005
R390 VSS.n31 VSS.t12 17.4005
R391 VSS.n31 VSS.t24 17.4005
R392 VSS.n57 VSS.n34 3.46248
R393 VSS.n50 VSS.n42 3.46248
R394 VSS.n48 VSS.n47 3.46248
R395 VSS.n41 VSS.n36 3.46248
R396 VSS.n93 VSS.n16 3.46248
R397 VSS.n89 VSS.n88 3.46248
R398 VSS.n101 VSS.n11 3.46248
R399 VSS.n98 VSS.n14 3.46248
R400 VSS.n106 VSS.n105 2.82278
R401 VSS.n4 VSS.n0 2.82278
R402 VSS.n111 VSS.n3 2.82278
R403 VSS.n74 VSS.n24 2.82278
R404 VSS.n72 VSS.n71 2.82278
R405 VSS.n70 VSS.n30 2.82278
R406 VSS.n59 VSS.n58 2.82278
R407 VSS.n102 VSS.n10 2.82278
R408 VSS.n49 VSS.n43 2.3255
R409 VSS.n56 VSS.n55 2.3255
R410 VSS.n100 VSS.n99 2.3255
R411 VSS.n92 VSS.n91 2.3255
R412 VSS.n73 VSS.n28 1.32907
R413 VSS.n69 VSS.n68 1.32907
R414 VSS.n113 VSS.n112 1.32907
R415 VSS.n104 VSS.n7 1.32907
R416 VSS.n24 VSS 0.90794
R417 VSS.n114 VSS.n2 0.685283
R418 VSS.n103 VSS.n9 0.685283
R419 VSS.n27 VSS.n26 0.685283
R420 VSS.n33 VSS.n32 0.685283
R421 VSS.n47 VSS 0.479667
R422 VSS VSS.n57 0.466646
R423 VSS VSS.n101 0.466646
R424 VSS.n71 VSS.n70 0.430188
R425 VSS.n105 VSS.n3 0.430188
R426 VSS.n89 VSS 0.404146
R427 VSS.n71 VSS.n28 0.359875
R428 VSS.n70 VSS.n69 0.359875
R429 VSS.n113 VSS.n3 0.359875
R430 VSS.n105 VSS.n104 0.359875
R431 VSS.n28 VSS.n27 0.229667
R432 VSS.n69 VSS.n33 0.229667
R433 VSS.n114 VSS.n113 0.229667
R434 VSS.n104 VSS.n103 0.229667
R435 VSS VSS.n0 0.191906
R436 VSS.n57 VSS.n56 0.189302
R437 VSS.n43 VSS.n42 0.189302
R438 VSS.n101 VSS.n100 0.189302
R439 VSS.n91 VSS.n16 0.189302
R440 VSS.n42 VSS.n41 0.141125
R441 VSS.n16 VSS.n14 0.141125
R442 VSS.n41 VSS.n35 0.13201
R443 VSS.n47 VSS.n46 0.13201
R444 VSS.n14 VSS.n12 0.13201
R445 VSS.n90 VSS.n89 0.13201
R446 VSS.n58 VSS.n33 0.130708
R447 VSS.n103 VSS.n102 0.130708
R448 VSS.n27 VSS 0.124198
R449 VSS VSS.n114 0.124198
R450 VSS.n58 VSS 0.0695104
R451 VSS.n102 VSS 0.0695104
R452 VSS.n56 VSS.n35 0.0577917
R453 VSS.n46 VSS.n43 0.0577917
R454 VSS.n100 VSS.n12 0.0577917
R455 VSS.n91 VSS.n90 0.0577917
R456 VSS VSS.n24 0.00701042
R457 VSS VSS.n0 0.00701042
R458 variable_delay_unit_1.forward.n0 variable_delay_unit_1.forward.t2 607.409
R459 variable_delay_unit_1.forward.n0 variable_delay_unit_1.forward.t3 321.423
R460 variable_delay_unit_1.forward variable_delay_unit_1.forward.n0 161.72
R461 variable_delay_unit_1.forward.n1 variable_delay_unit_1.forward.t1 84.7227
R462 variable_delay_unit_1.forward.n1 variable_delay_unit_1.forward.t0 84.0867
R463 variable_delay_unit_1.forward.n2 variable_delay_unit_1.forward 19.8934
R464 variable_delay_unit_1.forward variable_delay_unit_1.forward.n2 0.851271
R465 variable_delay_unit_1.forward.n2 variable_delay_unit_1.forward.n1 0.465495
R466 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t3 628.097
R467 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.t5 622.766
R468 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t7 523.774
R469 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t6 304.647
R470 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t2 304.647
R471 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t4 202.44
R472 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n0 168.969
R473 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n4 166.147
R474 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R475 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R476 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R477 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en 5.58443
R478 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n2 4.59003
R479 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.n3 1.09595
R480 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t2 607.409
R481 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t4 543.053
R482 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t3 321.423
R483 variable_delay_unit_1.in variable_delay_unit_1.in.n2 221.778
R484 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t5 221.72
R485 variable_delay_unit_1.in variable_delay_unit_1.in.n0 161.72
R486 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t0 84.7227
R487 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t1 84.0867
R488 variable_delay_unit_1.in.n3 variable_delay_unit_1.in 20.0791
R489 variable_delay_unit_1.in variable_delay_unit_1.in.n3 0.851271
R490 variable_delay_unit_1.in.n3 variable_delay_unit_1.in.n1 0.465495
R491 out.n0 out.t0 84.8477
R492 out.n2 out.t3 84.8477
R493 out.n0 out.t1 84.2063
R494 out.n2 out.t2 84.1683
R495 out out.n3 10.0241
R496 out.n1 out 0.681535
R497 out out.n0 0.287138
R498 out.n3 out 0.0803611
R499 out.n3 out.n2 0.0508472
R500 out.n1 out 0.013431
R501 out out.n1 0.0109167
R502 in.n0 in.t0 543.053
R503 in.n0 in.t1 221.72
R504 in in.n0 221.565
C0 VDD a_4562_352# 0.160518f
C1 variable_delay_unit_0.tristate_inverter_1.en a_1614_772# 0.11539f
C2 variable_delay_unit_1.tristate_inverter_1.en VDD 3.86972f
C3 VDD variable_delay_unit_1.out 1.61031f
C4 a_2496_352# a_2496_772# 0.011184f
C5 variable_delay_unit_1.tristate_inverter_1.en out 0.002141f
C6 out variable_delay_unit_1.out 0.071795f
C7 variable_delay_unit_1.forward a_4562_772# 0.088132f
C8 in variable_delay_unit_1.in 0.08442f
C9 variable_delay_unit_1.tristate_inverter_1.en a_5444_772# 0.029284f
C10 a_5444_772# variable_delay_unit_1.out 0.493816f
C11 variable_delay_unit_0.tristate_inverter_1.en a_2496_352# 0.15982f
C12 a_4562_352# variable_delay_unit_1.forward 0.054206f
C13 variable_delay_unit_1.out a_2496_772# 0.071074f
C14 variable_delay_unit_1.in a_1614_772# 0.088132f
C15 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.forward 0.794183f
C16 variable_delay_unit_1.forward variable_delay_unit_1.out 0.234428f
C17 VDD out 1.37861f
C18 in a_1614_772# 8.82e-20
C19 variable_delay_unit_1.in a_5444_352# 7.65e-21
C20 VDD a_5444_772# 1.78268f
C21 VDD a_1614_352# 0.160518f
C22 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en 0.002365f
C23 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.out 0.085059f
C24 VDD a_2496_772# 1.78275f
C25 out a_1614_352# 0.222585f
C26 VDD variable_delay_unit_1.forward 2.28565f
C27 out a_2496_772# 0.493816f
C28 a_4562_772# variable_delay_unit_1.in 8.82e-20
C29 in a_2496_352# 7.65e-21
C30 VDD variable_delay_unit_0.tristate_inverter_1.en 3.86872f
C31 a_4562_352# variable_delay_unit_1.in 8.82e-20
C32 a_5444_772# variable_delay_unit_1.forward 0.016896f
C33 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.in 0.09141f
C34 variable_delay_unit_0.tristate_inverter_1.en out 0.12022f
C35 variable_delay_unit_1.in variable_delay_unit_1.out 0.499092f
C36 variable_delay_unit_0.tristate_inverter_1.en a_1614_352# 2.39e-19
C37 variable_delay_unit_0.tristate_inverter_1.en a_2496_772# 0.029284f
C38 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.forward 7.91e-21
C39 VDD variable_delay_unit_1.in 3.20907f
C40 variable_delay_unit_1.tristate_inverter_1.en a_5444_352# 0.15982f
C41 variable_delay_unit_1.out a_5444_352# 0.172055f
C42 VDD in 0.498166f
C43 out variable_delay_unit_1.in 0.235655f
C44 out in 0.487038f
C45 VDD a_1614_772# 1.70112f
C46 a_5444_772# variable_delay_unit_1.in 7.65e-21
C47 a_1614_352# variable_delay_unit_1.in 0.054206f
C48 a_4562_352# a_4562_772# 0.004142f
C49 a_2496_352# variable_delay_unit_1.out 0.070146f
C50 VDD a_5444_352# 0.003377f
C51 in a_1614_352# 8.82e-20
C52 variable_delay_unit_1.in a_2496_772# 0.020173f
C53 variable_delay_unit_1.tristate_inverter_1.en a_4562_772# 0.11539f
C54 out a_1614_772# 0.505512f
C55 a_4562_772# variable_delay_unit_1.out 0.505512f
C56 variable_delay_unit_1.forward variable_delay_unit_1.in 0.087283f
C57 in a_2496_772# 7.65e-21
C58 variable_delay_unit_1.tristate_inverter_1.en a_4562_352# 2.39e-19
C59 a_4562_352# variable_delay_unit_1.out 0.222585f
C60 a_1614_352# a_1614_772# 0.004142f
C61 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.out 0.12029f
C62 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.in 0.814958f
C63 VDD a_2496_352# 0.003447f
C64 a_5444_772# a_5444_352# 0.011184f
C65 variable_delay_unit_0.tristate_inverter_1.en in 0.091118f
C66 VDD a_4562_772# 1.70112f
C67 out a_2496_352# 0.172055f
C68 out VSS 1.89289f
C69 in VSS 1.0591f
C70 VDD VSS 21.536554f
C71 a_5444_352# VSS 0.784074f
C72 a_4562_352# VSS 0.71648f
C73 a_2496_352# VSS 0.717347f
C74 a_1614_352# VSS 0.71648f
C75 a_5444_772# VSS 0.114203f
C76 a_4562_772# VSS 0.037888f
C77 variable_delay_unit_1.forward VSS 2.632682f
C78 variable_delay_unit_1.tristate_inverter_1.en VSS 2.962361f
C79 a_2496_772# VSS 0.043128f
C80 variable_delay_unit_1.out VSS 2.29732f
C81 a_1614_772# VSS 0.037888f
C82 variable_delay_unit_1.in VSS 4.167534f
C83 variable_delay_unit_0.tristate_inverter_1.en VSS 2.857091f
C84 variable_delay_unit_1.in.t2 VSS 0.068546f
C85 variable_delay_unit_1.in.t3 VSS 0.025993f
C86 variable_delay_unit_1.in.n0 VSS 0.072091f
C87 variable_delay_unit_1.in.t1 VSS 0.050497f
C88 variable_delay_unit_1.in.t0 VSS 0.160539f
C89 variable_delay_unit_1.in.n1 VSS 0.389091f
C90 variable_delay_unit_1.in.t4 VSS 0.065437f
C91 variable_delay_unit_1.in.t5 VSS 0.021123f
C92 variable_delay_unit_1.in.n2 VSS 0.068813f
C93 variable_delay_unit_1.in.n3 VSS 0.640809f
C94 variable_delay_unit_0.tristate_inverter_1.en.t4 VSS 0.027086f
C95 variable_delay_unit_0.tristate_inverter_1.en.t2 VSS 0.035f
C96 variable_delay_unit_0.tristate_inverter_1.en.t6 VSS 0.035f
C97 variable_delay_unit_0.tristate_inverter_1.en.n0 VSS 0.103163f
C98 variable_delay_unit_0.tristate_inverter_1.en.t1 VSS 0.215011f
C99 variable_delay_unit_0.tristate_inverter_1.en.t0 VSS 0.067642f
C100 variable_delay_unit_0.tristate_inverter_1.en.n1 VSS 0.85898f
C101 variable_delay_unit_0.tristate_inverter_1.en.n2 VSS 0.944443f
C102 variable_delay_unit_0.tristate_inverter_1.en.t5 VSS 0.093268f
C103 variable_delay_unit_0.tristate_inverter_1.en.t7 VSS 0.086397f
C104 variable_delay_unit_0.tristate_inverter_1.en.t3 VSS 0.093582f
C105 variable_delay_unit_0.tristate_inverter_1.en.n3 VSS 0.091588f
C106 variable_delay_unit_0.tristate_inverter_1.en.n4 VSS 0.06359f
C107 variable_delay_unit_1.forward.t2 VSS 0.067654f
C108 variable_delay_unit_1.forward.t3 VSS 0.025654f
C109 variable_delay_unit_1.forward.n0 VSS 0.071153f
C110 variable_delay_unit_1.forward.t0 VSS 0.04984f
C111 variable_delay_unit_1.forward.t1 VSS 0.15845f
C112 variable_delay_unit_1.forward.n1 VSS 0.384027f
C113 variable_delay_unit_1.forward.n2 VSS 0.632469f
C114 variable_delay_unit_1.tristate_inverter_1.en.t5 VSS 0.027086f
C115 variable_delay_unit_1.tristate_inverter_1.en.t2 VSS 0.035f
C116 variable_delay_unit_1.tristate_inverter_1.en.t3 VSS 0.035f
C117 variable_delay_unit_1.tristate_inverter_1.en.n0 VSS 0.103163f
C118 variable_delay_unit_1.tristate_inverter_1.en.t1 VSS 0.215011f
C119 variable_delay_unit_1.tristate_inverter_1.en.t0 VSS 0.067642f
C120 variable_delay_unit_1.tristate_inverter_1.en.n1 VSS 0.85898f
C121 variable_delay_unit_1.tristate_inverter_1.en.n2 VSS 0.944443f
C122 variable_delay_unit_1.tristate_inverter_1.en.t7 VSS 0.093268f
C123 variable_delay_unit_1.tristate_inverter_1.en.t4 VSS 0.086397f
C124 variable_delay_unit_1.tristate_inverter_1.en.t6 VSS 0.093582f
C125 variable_delay_unit_1.tristate_inverter_1.en.n3 VSS 0.091588f
C126 variable_delay_unit_1.tristate_inverter_1.en.n4 VSS 0.06359f
C127 VDD.n0 VSS 0.190382f
C128 VDD.t21 VSS 0.046888f
C129 VDD.n1 VSS 0.048588f
C130 VDD.n2 VSS 0.043398f
C131 VDD.n3 VSS 0.028635f
C132 VDD.t37 VSS 0.195867f
C133 VDD.n4 VSS 0.05654f
C134 VDD.n5 VSS 0.05654f
C135 VDD.t38 VSS 0.046888f
C136 VDD.n6 VSS 0.019547f
C137 VDD.n7 VSS 0.190382f
C138 VDD.n8 VSS 0.053221f
C139 VDD.t41 VSS 0.012494f
C140 VDD.t43 VSS 0.012494f
C141 VDD.n9 VSS 0.036465f
C142 VDD.t10 VSS 0.046131f
C143 VDD.n10 VSS 0.166326f
C144 VDD.n11 VSS 0.071912f
C145 VDD.n12 VSS 0.053221f
C146 VDD.n13 VSS 0.03368f
C147 VDD.n14 VSS 0.183676f
C148 VDD.t0 VSS 0.156929f
C149 VDD.n15 VSS 0.08687f
C150 VDD.n16 VSS 0.08687f
C151 VDD.t24 VSS 0.012494f
C152 VDD.t30 VSS 0.012494f
C153 VDD.n17 VSS 0.036465f
C154 VDD.t36 VSS 0.046131f
C155 VDD.n18 VSS 0.166326f
C156 VDD.t29 VSS 0.089287f
C157 VDD.n19 VSS 0.059525f
C158 VDD.t23 VSS 0.089287f
C159 VDD.t35 VSS 0.176037f
C160 VDD.n20 VSS 0.183676f
C161 VDD.n21 VSS 0.053345f
C162 VDD.n22 VSS 0.033479f
C163 VDD.n23 VSS 0.031158f
C164 VDD.n24 VSS 0.071912f
C165 VDD.n25 VSS 0.053221f
C166 VDD.n26 VSS 0.03368f
C167 VDD.n27 VSS 0.320623f
C168 VDD.n28 VSS 0.320623f
C169 VDD.t39 VSS 0.156929f
C170 VDD.t40 VSS 0.089287f
C171 VDD.t9 VSS 0.176037f
C172 VDD.t42 VSS 0.089287f
C173 VDD.n29 VSS 0.059525f
C174 VDD.n30 VSS 0.08687f
C175 VDD.n31 VSS 0.08687f
C176 VDD.n32 VSS 0.031158f
C177 VDD.n33 VSS 0.033824f
C178 VDD.n34 VSS 0.040685f
C179 VDD.n35 VSS 0.067617f
C180 VDD.n36 VSS 0.013029f
C181 VDD.n37 VSS 0.086505f
C182 VDD.n38 VSS 0.045555f
C183 VDD.n39 VSS 0.043398f
C184 VDD.n40 VSS 0.028635f
C185 VDD.n41 VSS 0.15551f
C186 VDD.n42 VSS 0.15551f
C187 VDD.t20 VSS 0.195867f
C188 VDD.n43 VSS 0.019547f
C189 VDD.n44 VSS 0.05654f
C190 VDD.n45 VSS 0.05654f
C191 VDD.n46 VSS 0.013029f
C192 VDD.n47 VSS 0.086505f
C193 VDD.n48 VSS 0.04795f
C194 VDD.t44 VSS 0.005903f
C195 VDD.t50 VSS 0.007627f
C196 VDD.t49 VSS 0.007627f
C197 VDD.n49 VSS 0.022481f
C198 VDD.t22 VSS 0.018828f
C199 VDD.t34 VSS 0.020394f
C200 VDD.n50 VSS 0.019959f
C201 VDD.t28 VSS 0.020325f
C202 VDD.n51 VSS 0.013858f
C203 VDD.n52 VSS 0.145601f
C204 VDD.n53 VSS 0.114252f
C205 VDD.t19 VSS 0.019086f
C206 VDD.t47 VSS 0.006161f
C207 VDD.n54 VSS 0.018816f
C208 VDD.n55 VSS 0.135399f
C209 VDD.n56 VSS 0.042655f
C210 VDD.n57 VSS 0.053221f
C211 VDD.t18 VSS 0.012494f
C212 VDD.t15 VSS 0.012494f
C213 VDD.n58 VSS 0.036465f
C214 VDD.t33 VSS 0.046131f
C215 VDD.n59 VSS 0.166326f
C216 VDD.n60 VSS 0.071912f
C217 VDD.n61 VSS 0.08687f
C218 VDD.n62 VSS 0.183676f
C219 VDD.t32 VSS 0.176037f
C220 VDD.t17 VSS 0.089287f
C221 VDD.n63 VSS 0.059525f
C222 VDD.t14 VSS 0.089287f
C223 VDD.t8 VSS 0.156929f
C224 VDD.t3 VSS 0.156929f
C225 VDD.n64 VSS 0.08687f
C226 VDD.n65 VSS 0.08687f
C227 VDD.t12 VSS 0.012494f
C228 VDD.t7 VSS 0.012494f
C229 VDD.n66 VSS 0.036465f
C230 VDD.t2 VSS 0.046131f
C231 VDD.n67 VSS 0.166326f
C232 VDD.t11 VSS 0.089287f
C233 VDD.n68 VSS 0.059525f
C234 VDD.t6 VSS 0.089287f
C235 VDD.t1 VSS 0.176037f
C236 VDD.n69 VSS 0.183676f
C237 VDD.n70 VSS 0.053221f
C238 VDD.n71 VSS 0.190382f
C239 VDD.t5 VSS 0.046888f
C240 VDD.n72 VSS 0.086505f
C241 VDD.n73 VSS 0.05654f
C242 VDD.n74 VSS 0.028635f
C243 VDD.n75 VSS 0.043398f
C244 VDD.t27 VSS 0.046888f
C245 VDD.n76 VSS 0.086505f
C246 VDD.n77 VSS 0.05654f
C247 VDD.t51 VSS 0.005903f
C248 VDD.t48 VSS 0.007627f
C249 VDD.t46 VSS 0.007627f
C250 VDD.n78 VSS 0.022481f
C251 VDD.t16 VSS 0.018828f
C252 VDD.t31 VSS 0.020394f
C253 VDD.n79 VSS 0.019959f
C254 VDD.t13 VSS 0.020325f
C255 VDD.n80 VSS 0.013858f
C256 VDD.n81 VSS 0.145601f
C257 VDD.n82 VSS 0.113749f
C258 VDD.t25 VSS 0.019086f
C259 VDD.t45 VSS 0.006161f
C260 VDD.n83 VSS 0.018825f
C261 VDD.n84 VSS 0.135893f
C262 VDD.n85 VSS 0.038385f
C263 VDD.n86 VSS 0.049068f
C264 VDD.n87 VSS 0.019547f
C265 VDD.t4 VSS 0.195867f
C266 VDD.n88 VSS 0.15551f
C267 VDD.n89 VSS 0.028635f
C268 VDD.n90 VSS 0.15551f
C269 VDD.t26 VSS 0.195867f
C270 VDD.n91 VSS 0.019547f
C271 VDD.n92 VSS 0.190382f
C272 VDD.n93 VSS 0.05654f
C273 VDD.n94 VSS 0.013029f
C274 VDD.n95 VSS 0.048588f
C275 VDD.n96 VSS 0.045555f
C276 VDD.n97 VSS 0.043398f
C277 VDD.n98 VSS 0.05654f
C278 VDD.n99 VSS 0.013029f
C279 VDD.n100 VSS 0.067617f
C280 VDD.n101 VSS 0.040685f
C281 VDD.n102 VSS 0.033824f
C282 VDD.n103 VSS 0.031158f
C283 VDD.n104 VSS 0.071912f
C284 VDD.n105 VSS 0.053221f
C285 VDD.n106 VSS 0.03368f
C286 VDD.n107 VSS 0.320623f
C287 VDD.n108 VSS 0.320623f
C288 VDD.n109 VSS 0.03368f
C289 VDD.n110 VSS 0.053221f
C290 VDD.n111 VSS 0.08687f
C291 VDD.n112 VSS 0.031158f
C292 VDD.n113 VSS 0.033479f
C293 VDD.n114 VSS 0.034136f
.ends

