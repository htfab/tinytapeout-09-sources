* NGSPICE file created from vernier_delay_line_parax.ext - technology: sky130A

.subckt vernier_delay_line_parax term_1 term_2 term_3 term_4 term_5 term_6 term_7
+ stop_strong start_neg start_pos VDD VSS term_0
X0 a_17348_1376# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VDD.t198 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 a_3116_2192.t5 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X2 VSS.t140 stop_strong.t0 a_11980_2192.t10 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X3 saff_delay_unit_5/delay_unit_2_0.in_1.t3 saff_delay_unit_4/delay_unit_2_0.in_2.t8 VSS.t369 VSS.t368 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X4 a_16632_2192# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X5 saff_delay_unit_3/delay_unit_2_0.in_2.t5 saff_delay_unit_2/delay_unit_2_0.in_1.t8 VDD.t178 VDD.t177 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X6 VSS.t308 start_pos.t2 start_neg.t0 VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X7 saff_delay_unit_2/delay_unit_2_0.in_1.t5 saff_delay_unit_1/delay_unit_2_0.in_2.t8 VSS.t319 VSS.t318 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X8 a_570_2192.t12 saff_delay_unit_1/delay_unit_2_0.in_2.t9 a_834_2192.t5 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X9 a_16544_2192.t12 saff_delay_unit_7/saff_2_0.d.t8 a_16632_2192# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X10 a_7804_296# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 term_3.t2 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 VDD.t71 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 a_14382_160# VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X12 a_14350_2192# saff_delay_unit_7/delay_unit_2_0.in_1.t8 a_14262_2192.t3 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X13 VSS.t142 stop_strong.t1 a_2852_2192.t8 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X14 a_570_2192.t11 saff_delay_unit_1/delay_unit_2_0.in_2.t10 a_834_2192.t4 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X15 VDD.t182 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 saff_delay_unit_3/saff_2_0.nq VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X16 term_7.t2 a_16664_160# VSS.t331 VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X17 saff_delay_unit_5/delay_unit_2_0.in_2.t2 saff_delay_unit_4/delay_unit_2_0.in_1.t8 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X18 a_3618_296# term_1.t4 VSS.t354 VSS.t353 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X19 VDD.t271 saff_delay_unit_7/saff_2_0.nq a_16932_730# VDD.t270 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X20 saff_delay_unit_4/delay_unit_2_0.in_2.t5 saff_delay_unit_3/delay_unit_2_0.in_1.t8 VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X21 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 a_16808_2192.t5 VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X22 saff_delay_unit_3/delay_unit_2_0.in_1.t4 saff_delay_unit_2/delay_unit_2_0.in_2.t8 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X23 VSS.t316 saff_delay_unit_1/delay_unit_2_0.in_2.t11 saff_delay_unit_1/delay_unit_2_0.in_1.t6 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X24 a_5398_2192.t4 saff_delay_unit_3/delay_unit_2_0.in_2.t8 a_5134_2192.t0 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X25 delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.d.t9 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X26 a_9786_2192# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X27 saff_delay_unit_7/saff_2_0.d.t3 saff_delay_unit_7/delay_unit_2_0.in_2.t8 VSS.t160 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X28 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X29 term_5.t1 a_12100_160# VSS.t187 VSS.t186 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X30 VSS.t27 saff_delay_unit_6/delay_unit_2_0.in_2.t8 saff_delay_unit_7/delay_unit_2_0.in_1.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X31 VSS.t385 stop_strong.t2 a_16544_2192.t8 VSS.t384 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X32 a_658_2192# saff_delay_unit_1/delay_unit_2_0.in_1.t8 a_570_2192.t2 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X33 a_5938_1376# saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X34 a_7804_730# a_7536_160# term_3.t1 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X35 a_7504_2192# saff_delay_unit_4/delay_unit_2_0.in_1.t9 a_7416_2192.t3 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X36 delay_unit_2_0.out_1.t5 saff_delay_unit_7/saff_2_0.nd.t8 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X37 VSS.t337 saff_delay_unit_6/delay_unit_2_0.in_1.t8 saff_delay_unit_7/delay_unit_2_0.in_2.t7 VSS.t336 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X38 a_17310_296# term_7.t4 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X39 VDD.t303 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VDD.t302 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X40 VDD.t115 saff_delay_unit_7/delay_unit_2_0.in_2.t9 saff_delay_unit_7/delay_unit_2_0.in_1.t4 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X41 saff_delay_unit_6/delay_unit_2_0.in_2.t3 saff_delay_unit_5/delay_unit_2_0.in_1.t8 VSS.t246 VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X42 a_7504_2192# saff_delay_unit_4/delay_unit_2_0.in_1.t10 a_7416_2192.t2 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X43 VDD.t202 start_neg.t2 saff_delay_unit_1/delay_unit_2_0.in_1.t5 VDD.t201 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X44 term_7.t1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X45 VSS.t227 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 a_2972_160# VSS.t226 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X46 a_12068_2192# saff_delay_unit_6/delay_unit_2_0.in_1.t9 a_11980_2192.t4 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X47 a_3618_730# term_1.t5 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X48 a_9698_2192.t12 saff_delay_unit_5/delay_unit_2_0.in_2.t8 a_9962_2192.t0 VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X49 saff_delay_unit_7/delay_unit_2_0.in_2.t5 saff_delay_unit_6/delay_unit_2_0.in_1.t10 VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X50 VSS.t387 stop_strong.t3 a_11980_2192.t9 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X51 VSS.t25 saff_delay_unit_7/delay_unit_2_0.in_1.t9 saff_delay_unit_7/delay_unit_2_0.in_2.t1 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X52 saff_delay_unit_6/delay_unit_2_0.in_1.t4 saff_delay_unit_5/delay_unit_2_0.in_2.t9 VSS.t232 VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X53 VDD.t81 saff_delay_unit_1/delay_unit_2_0.in_1.t9 saff_delay_unit_1/delay_unit_2_0.in_2.t1 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X54 saff_delay_unit_2/saff_2_0.nq saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 a_5900_296# VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X55 VSS.t74 saff_delay_unit_2/saff_2_0.nq a_5522_296# VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X56 VSS.t295 saff_delay_unit_3/delay_unit_2_0.in_2.t9 saff_delay_unit_4/delay_unit_2_0.in_1.t2 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X57 VSS.t310 start_pos.t3 saff_delay_unit_1/delay_unit_2_0.in_2.t4 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X58 term_5.t0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X59 term_0.t1 a_690_160# VSS.t71 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X60 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 a_14350_2192# VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X61 VDD.t313 saff_delay_unit_5/delay_unit_2_0.in_2.t10 saff_delay_unit_5/delay_unit_2_0.in_1.t7 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X62 a_2940_2192# saff_delay_unit_2/delay_unit_2_0.in_1.t9 a_2852_2192.t12 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X63 VSS.t37 stop_strong.t4 a_2852_2192.t7 VSS.t36 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X64 a_5938_1376# saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X65 a_14526_2192.t5 saff_delay_unit_7/delay_unit_2_0.in_2.t10 a_14262_2192.t7 VSS.t178 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X66 a_570_2192.t8 stop_strong.t5 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X67 saff_delay_unit_3/delay_unit_2_0.in_2.t2 saff_delay_unit_2/delay_unit_2_0.in_1.t10 VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X68 a_14650_296# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 term_6.t0 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X69 a_17310_730# term_7.t5 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X70 a_11980_2192.t2 saff_delay_unit_6/delay_unit_2_0.in_1.t11 a_12068_2192# VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X71 VDD.t65 saff_delay_unit_4/delay_unit_2_0.in_2.t9 saff_delay_unit_4/delay_unit_2_0.in_1.t7 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X72 saff_delay_unit_0/saff_2_0.nq saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 a_1336_296# VSS.t340 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X73 a_14526_2192.t4 saff_delay_unit_7/delay_unit_2_0.in_2.t11 a_14262_2192.t4 VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X74 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 stop_strong.t6 VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X75 saff_delay_unit_7/saff_2_0.nd.t2 saff_delay_unit_7/delay_unit_2_0.in_1.t10 VSS.t389 VSS.t388 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X76 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 a_5398_2192.t5 VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X77 VDD.t63 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 a_2972_160# VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X78 a_2852_2192.t2 saff_delay_unit_2/delay_unit_2_0.in_2.t9 a_3116_2192.t2 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X79 a_10464_296# term_4.t4 VSS.t205 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X80 saff_delay_unit_4/delay_unit_2_0.in_2.t0 saff_delay_unit_3/delay_unit_2_0.in_1.t9 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X81 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 a_9962_2192.t5 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X82 VSS.t220 stop_strong.t7 a_5134_2192.t8 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X83 a_2852_2192.t3 saff_delay_unit_2/delay_unit_2_0.in_2.t10 a_3116_2192.t3 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X84 term_2.t2 a_5254_160# VSS.t289 VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X85 VSS.t321 saff_delay_unit_1/delay_unit_2_0.in_2.t12 saff_delay_unit_2/delay_unit_2_0.in_1.t6 VSS.t320 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X86 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X87 VSS.t287 saff_delay_unit_4/delay_unit_2_0.in_1.t11 saff_delay_unit_4/delay_unit_2_0.in_2.t6 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X88 saff_delay_unit_2/saff_2_0.nq a_5938_1376# a_5900_730# VDD.t159 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X89 VSS.t362 stop_strong.t8 a_16544_2192.t7 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X90 a_16632_2192# saff_delay_unit_7/saff_2_0.d.t10 a_16544_2192.t11 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X91 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 a_7680_2192.t1 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X92 VDD.t47 saff_delay_unit_2/saff_2_0.nq a_5522_730# VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X93 term_0.t3 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X94 a_14262_2192.t12 stop_strong.t9 VSS.t364 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X95 a_12784_1376# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 VSS.t339 VSS.t338 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X96 delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.d.t11 VSS.t283 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X97 a_834_2192.t3 saff_delay_unit_1/delay_unit_2_0.in_2.t13 a_570_2192.t10 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X98 VDD.t15 saff_delay_unit_2/delay_unit_2_0.in_2.t11 saff_delay_unit_2/delay_unit_2_0.in_1.t1 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X99 VDD.t289 saff_delay_unit_7/delay_unit_2_0.in_2.t12 saff_delay_unit_7/saff_2_0.d.t5 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X100 saff_delay_unit_6/delay_unit_2_0.in_2.t2 saff_delay_unit_5/delay_unit_2_0.in_1.t9 VSS.t268 VSS.t267 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X101 a_14650_730# a_14382_160# term_6.t3 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X102 a_7680_2192.t5 saff_delay_unit_4/delay_unit_2_0.in_2.t10 a_7416_2192.t12 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X103 saff_delay_unit_7/delay_unit_2_0.in_1.t6 saff_delay_unit_6/delay_unit_2_0.in_2.t9 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X104 VSS.t391 saff_delay_unit_4/delay_unit_2_0.in_1.t12 saff_delay_unit_5/delay_unit_2_0.in_2.t1 VSS.t390 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X105 a_10086_296# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 term_4.t3 VSS.t173 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X106 a_5134_2192.t7 stop_strong.t10 VSS.t242 VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X107 saff_delay_unit_0/saff_2_0.nq a_1374_1376# a_1336_730# VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X108 saff_delay_unit_7/delay_unit_2_0.in_2.t6 saff_delay_unit_6/delay_unit_2_0.in_1.t12 VDD.t258 VDD.t257 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X109 saff_delay_unit_6/saff_2_0.nq saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 a_15028_296# VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X110 a_9698_2192.t3 saff_delay_unit_5/delay_unit_2_0.in_1.t10 a_9786_2192# VSS.t374 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X111 delay_unit_2_0.out_1.t2 saff_delay_unit_7/saff_2_0.nd.t9 VSS.t380 VSS.t379 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X112 VDD.t283 saff_delay_unit_5/delay_unit_2_0.in_1.t11 saff_delay_unit_5/delay_unit_2_0.in_2.t7 VDD.t282 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X113 a_16544_2192.t2 saff_delay_unit_7/saff_2_0.nd.t10 a_16808_2192.t2 VSS.t180 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X114 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X115 saff_delay_unit_3/delay_unit_2_0.in_1.t5 saff_delay_unit_2/delay_unit_2_0.in_2.t12 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X116 VSS.t91 a_3656_1376# saff_delay_unit_1/saff_2_0.nq VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X117 VSS.t291 start_neg.t3 start_pos.t1 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X118 a_10464_730# term_4.t5 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X119 a_834_2192.t0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X120 a_9698_2192.t8 stop_strong.t11 VSS.t244 VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X121 VSS.t395 saff_delay_unit_3/delay_unit_2_0.in_2.t10 saff_delay_unit_3/delay_unit_2_0.in_1.t6 VSS.t394 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X122 term_2.t1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VDD.t206 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X123 a_9786_2192# saff_delay_unit_5/delay_unit_2_0.in_1.t12 a_9698_2192.t2 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X124 VSS.t223 saff_delay_unit_7/delay_unit_2_0.in_1.t11 saff_delay_unit_7/saff_2_0.nd.t1 VSS.t222 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X125 VSS.t177 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 a_9818_160# VSS.t176 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X126 VDD.t79 saff_delay_unit_1/delay_unit_2_0.in_1.t10 saff_delay_unit_2/delay_unit_2_0.in_2.t5 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X127 VDD.t89 saff_delay_unit_7/saff_2_0.nd.t11 saff_delay_unit_7/saff_2_0.d.t2 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X128 saff_delay_unit_5/saff_2_0.nq saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 a_12746_296# VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X129 a_7416_2192.t8 stop_strong.t12 VSS.t342 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X130 VDD.t279 stop_strong.t13 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X131 a_12784_1376# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X132 VDD.t232 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VDD.t231 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X133 VDD.t132 saff_delay_unit_5/delay_unit_2_0.in_2.t11 saff_delay_unit_6/delay_unit_2_0.in_1.t7 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X134 a_570_2192.t7 stop_strong.t14 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X135 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 stop_strong.t15 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X136 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 a_5222_2192# VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X137 a_14350_2192# saff_delay_unit_7/delay_unit_2_0.in_1.t12 a_14262_2192.t2 VSS.t376 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X138 saff_delay_unit_3/delay_unit_2_0.in_2.t1 saff_delay_unit_2/delay_unit_2_0.in_1.t11 VSS.t124 VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X139 a_11980_2192.t1 saff_delay_unit_6/delay_unit_2_0.in_2.t10 a_12244_2192.t5 VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X140 VDD.t25 saff_delay_unit_4/delay_unit_2_0.in_2.t11 saff_delay_unit_5/delay_unit_2_0.in_1.t6 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X141 a_10086_730# a_9818_160# term_4.t1 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X142 VDD.t87 saff_delay_unit_2/delay_unit_2_0.in_1.t12 saff_delay_unit_2/delay_unit_2_0.in_2.t7 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X143 a_3240_296# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 term_1.t2 VSS.t259 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X144 VSS.t195 saff_delay_unit_5/saff_2_0.nq a_12368_296# VSS.t194 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X145 saff_delay_unit_6/saff_2_0.nq a_15066_1376# a_15028_730# VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X146 VDD.t105 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 saff_delay_unit_1/saff_2_0.nq VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X147 a_2852_2192.t11 saff_delay_unit_2/delay_unit_2_0.in_1.t13 a_2940_2192# VSS.t117 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X148 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X149 VDD.t29 saff_delay_unit_6/delay_unit_2_0.in_2.t11 saff_delay_unit_6/delay_unit_2_0.in_1.t1 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X150 saff_delay_unit_3/saff_2_0.nq saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 a_8182_296# VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X151 a_16808_2192.t1 saff_delay_unit_7/saff_2_0.nd.t12 a_16544_2192.t1 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X152 VSS.t261 a_17348_1376# saff_delay_unit_7/saff_2_0.nq VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X153 a_2852_2192.t6 stop_strong.t16 VSS.t254 VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X154 saff_delay_unit_4/delay_unit_2_0.in_2.t2 saff_delay_unit_3/delay_unit_2_0.in_1.t10 VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X155 VDD.t91 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 a_9818_160# VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X156 a_14262_2192.t11 stop_strong.t17 VSS.t256 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X157 a_14262_2192.t1 saff_delay_unit_7/delay_unit_2_0.in_1.t13 a_14350_2192# VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X158 saff_delay_unit_5/saff_2_0.nq a_12784_1376# a_12746_730# VDD.t221 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X159 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 stop_strong.t18 VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X160 VDD.t1 saff_delay_unit_2/delay_unit_2_0.in_2.t13 saff_delay_unit_3/delay_unit_2_0.in_1.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X161 saff_delay_unit_2/delay_unit_2_0.in_1.t7 saff_delay_unit_1/delay_unit_2_0.in_2.t14 VDD.t252 VDD.t251 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X162 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 stop_strong.t19 VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X163 delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.d.t12 VSS.t266 VSS.t265 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X164 a_5134_2192.t3 saff_delay_unit_3/delay_unit_2_0.in_2.t11 a_5398_2192.t3 VSS.t396 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X165 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 a_12244_2192.t1 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X166 VDD.t130 saff_delay_unit_7/saff_2_0.d.t13 saff_delay_unit_7/saff_2_0.nd.t7 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X167 saff_delay_unit_7/delay_unit_2_0.in_1.t2 saff_delay_unit_6/delay_unit_2_0.in_2.t12 VDD.t57 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X168 a_1374_1376# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X169 a_5134_2192.t1 saff_delay_unit_3/delay_unit_2_0.in_2.t12 a_5398_2192.t2 VSS.t348 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X170 delay_unit_2_0.out_1.t1 saff_delay_unit_7/saff_2_0.nd.t13 VSS.t273 VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X171 a_16544_2192.t10 saff_delay_unit_7/saff_2_0.d.t14 a_16632_2192# VSS.t228 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X172 VDD.t297 saff_delay_unit_5/delay_unit_2_0.in_1.t13 saff_delay_unit_6/delay_unit_2_0.in_2.t6 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X173 VSS.t81 saff_delay_unit_7/delay_unit_2_0.in_2.t13 saff_delay_unit_7/delay_unit_2_0.in_1.t1 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X174 a_3240_730# a_2972_160# term_1.t1 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X175 saff_delay_unit_5/delay_unit_2_0.in_2.t5 saff_delay_unit_4/delay_unit_2_0.in_1.t13 VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X176 VDD.t163 saff_delay_unit_5/saff_2_0.nq a_12368_730# VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X177 a_9698_2192.t11 saff_delay_unit_5/delay_unit_2_0.in_2.t12 a_9962_2192.t2 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X178 a_7680_2192.t0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X179 VSS.t293 start_neg.t4 saff_delay_unit_1/delay_unit_2_0.in_1.t2 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X180 VSS.t153 a_10502_1376# saff_delay_unit_4/saff_2_0.nq VSS.t152 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X181 a_9698_2192.t7 stop_strong.t20 VSS.t216 VSS.t215 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X182 a_7416_2192.t9 saff_delay_unit_4/delay_unit_2_0.in_2.t12 a_7680_2192.t4 VSS.t99 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X183 saff_delay_unit_3/saff_2_0.nq a_8220_1376# a_8182_730# VDD.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X184 a_12068_2192# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X185 VDD.t256 saff_delay_unit_7/saff_2_0.nd.t14 delay_unit_2_0.out_1.t4 VDD.t255 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X186 saff_delay_unit_7/delay_unit_2_0.in_2.t0 saff_delay_unit_6/delay_unit_2_0.in_1.t13 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X187 VDD.t234 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 saff_delay_unit_7/saff_2_0.nq VDD.t233 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X188 a_9962_2192.t1 saff_delay_unit_5/delay_unit_2_0.in_2.t13 a_9698_2192.t10 VSS.t269 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X189 saff_delay_unit_1/delay_unit_2_0.in_2.t7 start_pos.t4 VDD.t242 VDD.t241 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X190 saff_delay_unit_7/saff_2_0.d.t1 saff_delay_unit_7/delay_unit_2_0.in_2.t14 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X191 a_7416_2192.t7 stop_strong.t21 VSS.t218 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X192 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 stop_strong.t22 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X193 VSS.t113 saff_delay_unit_1/delay_unit_2_0.in_1.t11 saff_delay_unit_1/delay_unit_2_0.in_2.t0 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X194 saff_delay_unit_7/saff_2_0.nd.t5 saff_delay_unit_7/delay_unit_2_0.in_1.t14 VDD.t187 VDD.t186 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X195 VDD.t43 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X196 term_3.t0 a_7536_160# VSS.t189 VSS.t188 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X197 a_11980_2192.t5 saff_delay_unit_6/delay_unit_2_0.in_1.t14 a_12068_2192# VSS.t196 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X198 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X199 VSS.t240 saff_delay_unit_5/delay_unit_2_0.in_2.t14 saff_delay_unit_5/delay_unit_2_0.in_1.t0 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X200 saff_delay_unit_4/delay_unit_2_0.in_1.t5 saff_delay_unit_3/delay_unit_2_0.in_2.t13 VDD.t317 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X201 a_9786_2192# saff_delay_unit_5/delay_unit_2_0.in_1.t14 a_9698_2192.t1 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X202 a_1374_1376# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X203 a_3116_2192.t4 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X204 VSS.t366 saff_delay_unit_4/delay_unit_2_0.in_2.t13 saff_delay_unit_4/delay_unit_2_0.in_1.t6 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X205 VSS.t304 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 a_16664_160# VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X206 VDD.t85 saff_delay_unit_2/delay_unit_2_0.in_1.t14 saff_delay_unit_3/delay_unit_2_0.in_2.t4 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X207 a_15066_1376# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VSS.t325 VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X208 a_834_2192.t2 saff_delay_unit_1/delay_unit_2_0.in_2.t15 a_570_2192.t9 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X209 VDD.t136 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 saff_delay_unit_4/saff_2_0.nq VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X210 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 a_658_2192# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X211 VDD.t109 stop_strong.t23 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X212 a_2852_2192.t5 stop_strong.t24 VSS.t149 VSS.t148 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X213 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 stop_strong.t25 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X214 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 a_7504_2192# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X215 VSS.t183 stop_strong.t26 a_570_2192.t6 VSS.t182 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X216 a_16632_2192# saff_delay_unit_7/saff_2_0.d.t15 a_16544_2192.t9 VSS.t184 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X217 VSS.t371 saff_delay_unit_0/saff_2_0.nq a_958_296# VSS.t370 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X218 saff_delay_unit_4/delay_unit_2_0.in_2.t4 saff_delay_unit_3/delay_unit_2_0.in_1.t11 VSS.t248 VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X219 VSS.t202 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 a_12100_160# VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X220 a_5134_2192.t12 saff_delay_unit_3/delay_unit_2_0.in_1.t12 a_5222_2192# VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X221 VSS.t191 a_5938_1376# saff_delay_unit_2/saff_2_0.nq VSS.t190 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X222 VDD.t200 saff_delay_unit_3/delay_unit_2_0.in_1.t13 saff_delay_unit_3/delay_unit_2_0.in_2.t6 VDD.t199 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X223 term_3.t3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VDD.t254 VDD.t253 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X224 a_5134_2192.t11 saff_delay_unit_3/delay_unit_2_0.in_1.t14 a_5222_2192# VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X225 a_5900_296# term_2.t4 VSS.t132 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X226 VSS.t1 saff_delay_unit_2/delay_unit_2_0.in_2.t14 saff_delay_unit_2/delay_unit_2_0.in_1.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X227 VDD.t69 saff_delay_unit_7/saff_2_0.d.t16 delay_unit_2_0.out_2 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X228 VSS.t378 saff_delay_unit_7/delay_unit_2_0.in_2.t15 saff_delay_unit_7/saff_2_0.d.t7 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X229 VDD.t152 stop_strong.t27 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VDD.t151 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X230 saff_delay_unit_7/delay_unit_2_0.in_1.t7 saff_delay_unit_6/delay_unit_2_0.in_2.t13 VSS.t347 VSS.t346 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X231 VDD.t236 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 a_16664_160# VDD.t235 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X232 a_15066_1376# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VDD.t277 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X233 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 a_2940_2192# VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X234 saff_delay_unit_7/delay_unit_2_0.in_2.t3 saff_delay_unit_6/delay_unit_2_0.in_1.t15 VSS.t95 VSS.t94 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X235 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 stop_strong.t28 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X236 VSS.t373 saff_delay_unit_5/delay_unit_2_0.in_1.t15 saff_delay_unit_5/delay_unit_2_0.in_2.t6 VSS.t372 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X237 saff_delay_unit_3/delay_unit_2_0.in_1.t1 saff_delay_unit_2/delay_unit_2_0.in_2.t15 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X238 VDD.t295 saff_delay_unit_0/saff_2_0.nq a_958_730# VDD.t294 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X239 a_7416_2192.t11 saff_delay_unit_4/delay_unit_2_0.in_2.t14 a_7680_2192.t3 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X240 a_5522_296# saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 term_2.t0 VSS.t158 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X241 saff_delay_unit_1/delay_unit_2_0.in_1.t4 start_neg.t5 VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X242 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 a_14526_2192.t1 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X243 VSS.t130 stop_strong.t29 a_5134_2192.t6 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X244 VDD.t41 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 a_12100_160# VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X245 VSS.t344 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 a_690_160# VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X246 VSS.t111 saff_delay_unit_1/delay_unit_2_0.in_1.t12 saff_delay_unit_2/delay_unit_2_0.in_2.t4 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X247 saff_delay_unit_4/delay_unit_2_0.in_1.t4 saff_delay_unit_3/delay_unit_2_0.in_2.t14 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X248 VDD.t95 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 saff_delay_unit_2/saff_2_0.nq VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X249 VSS.t41 saff_delay_unit_7/saff_2_0.nd.t15 saff_delay_unit_7/saff_2_0.d.t0 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X250 saff_delay_unit_1/delay_unit_2_0.in_2.t6 start_pos.t5 VDD.t244 VDD.t243 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X251 a_11980_2192.t11 saff_delay_unit_6/delay_unit_2_0.in_2.t14 a_12244_2192.t4 VSS.t271 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X252 term_6.t2 a_14382_160# VSS.t235 VSS.t234 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X253 VSS.t230 saff_delay_unit_5/delay_unit_2_0.in_2.t15 saff_delay_unit_6/delay_unit_2_0.in_1.t3 VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X254 a_5900_730# term_2.t5 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X255 a_8220_1376# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VSS.t210 VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X256 VSS.t98 saff_delay_unit_4/delay_unit_2_0.in_2.t15 saff_delay_unit_5/delay_unit_2_0.in_1.t2 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X257 a_7680_2192.t2 saff_delay_unit_4/delay_unit_2_0.in_2.t16 a_7416_2192.t10 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X258 saff_delay_unit_2/delay_unit_2_0.in_2.t3 saff_delay_unit_1/delay_unit_2_0.in_1.t13 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X259 VSS.t275 stop_strong.t30 a_570_2192.t5 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X260 VSS.t122 saff_delay_unit_2/delay_unit_2_0.in_1.t15 saff_delay_unit_2/delay_unit_2_0.in_2.t6 VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X261 a_12068_2192# saff_delay_unit_6/delay_unit_2_0.in_1.t16 a_11980_2192.t0 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X262 VDD.t180 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X263 VSS.t250 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 a_5254_160# VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X264 a_658_2192# saff_delay_unit_1/delay_unit_2_0.in_1.t14 a_570_2192.t3 VSS.t192 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X265 VSS.t48 saff_delay_unit_6/delay_unit_2_0.in_2.t15 saff_delay_unit_6/delay_unit_2_0.in_1.t0 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X266 saff_delay_unit_5/delay_unit_2_0.in_1.t5 saff_delay_unit_4/delay_unit_2_0.in_2.t17 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X267 a_5522_730# a_5254_160# term_2.t3 VDD.t224 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X268 VDD.t293 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 a_690_160# VDD.t292 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X269 VSS.t281 a_12784_1376# saff_delay_unit_5/saff_2_0.nq VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X270 a_3116_2192.t0 saff_delay_unit_2/delay_unit_2_0.in_2.t16 a_2852_2192.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X271 VDD.t189 saff_delay_unit_3/delay_unit_2_0.in_1.t15 saff_delay_unit_4/delay_unit_2_0.in_2.t3 VDD.t188 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X272 VSS.t333 saff_delay_unit_3/saff_2_0.nq a_7804_296# VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X273 a_9962_2192.t4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X274 VSS.t6 saff_delay_unit_2/delay_unit_2_0.in_2.t17 saff_delay_unit_3/delay_unit_2_0.in_1.t2 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X275 term_6.t1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 VDD.t165 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X276 a_3116_2192.t1 saff_delay_unit_2/delay_unit_2_0.in_2.t18 a_2852_2192.t1 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X277 saff_delay_unit_2/delay_unit_2_0.in_1.t2 saff_delay_unit_1/delay_unit_2_0.in_2.t16 VSS.t252 VSS.t251 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X278 VDD.t214 stop_strong.t31 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VDD.t213 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X279 a_8220_1376# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X280 a_16544_2192.t6 stop_strong.t32 VSS.t358 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X281 VSS.t360 stop_strong.t33 a_14262_2192.t10 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X282 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 a_9786_2192# VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X283 VDD.t21 stop_strong.t34 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X284 a_16932_296# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 term_7.t0 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X285 VSS.t77 saff_delay_unit_7/saff_2_0.d.t17 saff_delay_unit_7/saff_2_0.nd.t6 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X286 saff_delay_unit_7/delay_unit_2_0.in_1.t5 saff_delay_unit_6/delay_unit_2_0.in_2.t16 VSS.t157 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X287 a_570_2192.t1 saff_delay_unit_1/delay_unit_2_0.in_1.t15 a_658_2192# VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X288 saff_delay_unit_1/saff_2_0.nq saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 a_3618_296# VSS.t224 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X289 VSS.t45 saff_delay_unit_5/delay_unit_2_0.in_1.t16 saff_delay_unit_6/delay_unit_2_0.in_2.t1 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X290 VDD.t23 stop_strong.t35 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X291 a_7416_2192.t1 saff_delay_unit_4/delay_unit_2_0.in_1.t14 a_7504_2192# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X292 saff_delay_unit_5/delay_unit_2_0.in_2.t0 saff_delay_unit_4/delay_unit_2_0.in_1.t15 VSS.t208 VSS.t207 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X293 VSS.t87 stop_strong.t36 a_5134_2192.t5 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X294 VDD.t230 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 a_5254_160# VDD.t229 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X295 a_7416_2192.t0 saff_delay_unit_4/delay_unit_2_0.in_1.t16 a_7504_2192# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X296 a_12746_296# term_5.t4 VSS.t323 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X297 VDD.t307 saff_delay_unit_6/delay_unit_2_0.in_1.t17 saff_delay_unit_6/delay_unit_2_0.in_2.t7 VDD.t306 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X298 saff_delay_unit_1/delay_unit_2_0.in_1.t3 start_neg.t6 VDD.t275 VDD.t274 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X299 VDD.t39 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_5/saff_2_0.nq VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X300 VSS.t29 saff_delay_unit_7/saff_2_0.nd.t16 delay_unit_2_0.out_1.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X301 saff_delay_unit_1/delay_unit_2_0.in_2.t3 start_pos.t6 VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X302 saff_delay_unit_7/saff_2_0.d.t4 saff_delay_unit_7/delay_unit_2_0.in_2.t16 VSS.t214 VSS.t213 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X303 VDD.t267 saff_delay_unit_3/saff_2_0.nq a_7804_730# VDD.t266 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X304 VSS.t277 saff_delay_unit_1/saff_2_0.nq a_3240_296# VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X305 a_11980_2192.t8 stop_strong.t37 VSS.t89 VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X306 saff_delay_unit_7/saff_2_0.nd.t0 saff_delay_unit_7/delay_unit_2_0.in_1.t15 VSS.t352 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X307 saff_delay_unit_2/delay_unit_2_0.in_2.t2 saff_delay_unit_1/delay_unit_2_0.in_1.t16 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X308 VSS.t58 stop_strong.t38 a_7416_2192.t6 VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X309 a_2852_2192.t10 saff_delay_unit_2/delay_unit_2_0.in_1.t16 a_2940_2192# VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X310 saff_delay_unit_4/delay_unit_2_0.in_1.t1 saff_delay_unit_3/delay_unit_2_0.in_2.t15 VSS.t116 VSS.t115 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X311 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X312 a_16932_730# a_16664_160# term_7.t3 VDD.t265 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X313 term_1.t0 a_2972_160# VSS.t79 VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X314 a_12368_296# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 term_5.t3 VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X315 saff_delay_unit_6/delay_unit_2_0.in_1.t6 saff_delay_unit_5/delay_unit_2_0.in_2.t16 VDD.t285 VDD.t284 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X316 saff_delay_unit_1/saff_2_0.nq a_3656_1376# a_3618_730# VDD.t53 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X317 a_5222_2192# saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X318 a_14262_2192.t5 saff_delay_unit_7/delay_unit_2_0.in_2.t17 a_14526_2192.t3 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X319 VSS.t120 saff_delay_unit_2/delay_unit_2_0.in_1.t17 saff_delay_unit_3/delay_unit_2_0.in_2.t0 VSS.t119 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X320 a_12244_2192.t3 saff_delay_unit_6/delay_unit_2_0.in_2.t17 a_11980_2192.t3 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X321 saff_delay_unit_5/delay_unit_2_0.in_1.t4 saff_delay_unit_4/delay_unit_2_0.in_2.t18 VDD.t176 VDD.t175 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X322 VSS.t60 stop_strong.t39 a_11980_2192.t7 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X323 a_8182_296# term_3.t4 VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X324 saff_delay_unit_7/saff_2_0.nq saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 a_17310_296# VSS.t306 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X325 VDD.t240 start_pos.t7 start_neg.t1 VDD.t239 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X326 a_14262_2192.t6 saff_delay_unit_7/delay_unit_2_0.in_2.t18 a_14526_2192.t2 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X327 saff_delay_unit_2/delay_unit_2_0.in_1.t4 saff_delay_unit_1/delay_unit_2_0.in_2.t17 VDD.t248 VDD.t247 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X328 a_12746_730# term_5.t5 VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X329 VDD.t210 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X330 a_16808_2192.t4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X331 a_2940_2192# saff_delay_unit_2/delay_unit_2_0.in_1.t18 a_2852_2192.t9 VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X332 a_5134_2192.t4 stop_strong.t40 VSS.t83 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X333 VDD.t216 saff_delay_unit_1/saff_2_0.nq a_3240_730# VDD.t215 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X334 VSS.t85 stop_strong.t41 a_2852_2192.t4 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X335 VSS.t69 a_1374_1376# saff_delay_unit_0/saff_2_0.nq VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X336 a_10502_1376# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X337 saff_delay_unit_5/delay_unit_2_0.in_2.t4 saff_delay_unit_4/delay_unit_2_0.in_1.t17 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X338 VSS.t350 saff_delay_unit_3/delay_unit_2_0.in_1.t16 saff_delay_unit_3/delay_unit_2_0.in_2.t7 VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X339 a_16544_2192.t5 stop_strong.t42 VSS.t54 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X340 saff_delay_unit_3/delay_unit_2_0.in_1.t3 saff_delay_unit_2/delay_unit_2_0.in_2.t19 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X341 VSS.t56 stop_strong.t43 a_14262_2192.t9 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X342 term_1.t3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X343 a_12368_730# a_12100_160# term_5.t2 VDD.t157 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X344 VSS.t155 saff_delay_unit_7/saff_2_0.d.t18 delay_unit_2_0.out_2 VSS.t154 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X345 VDD.t250 saff_delay_unit_1/delay_unit_2_0.in_2.t18 saff_delay_unit_1/delay_unit_2_0.in_1.t7 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X346 a_958_296# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 term_0.t0 VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X347 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 a_10464_296# VSS.t355 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X348 a_5398_2192.t1 saff_delay_unit_3/delay_unit_2_0.in_2.t16 a_5134_2192.t2 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X349 saff_delay_unit_7/saff_2_0.d.t6 saff_delay_unit_7/delay_unit_2_0.in_2.t19 VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X350 a_8182_730# term_3.t5 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X351 VDD.t99 saff_delay_unit_6/delay_unit_2_0.in_2.t18 saff_delay_unit_7/delay_unit_2_0.in_1.t3 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X352 saff_delay_unit_7/saff_2_0.nq a_17348_1376# a_17310_730# VDD.t192 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X353 a_12244_2192.t0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X354 VSS.t279 saff_delay_unit_6/saff_2_0.nq a_14650_296# VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X355 VDD.t101 saff_delay_unit_6/delay_unit_2_0.in_1.t18 saff_delay_unit_7/delay_unit_2_0.in_2.t4 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X356 a_9962_2192.t3 saff_delay_unit_5/delay_unit_2_0.in_2.t17 a_9698_2192.t9 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X357 saff_delay_unit_6/delay_unit_2_0.in_2.t5 saff_delay_unit_5/delay_unit_2_0.in_1.t17 VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X358 VSS.t393 stop_strong.t44 a_16544_2192.t4 VSS.t392 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X359 VDD.t311 stop_strong.t45 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X360 saff_delay_unit_1/delay_unit_2_0.in_1.t1 start_neg.t7 VSS.t302 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X361 VSS.t285 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 a_7536_160# VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X362 a_1336_296# term_0.t4 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X363 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 a_834_2192.t1 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X364 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 a_16632_2192# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X365 VSS.t136 stop_strong.t46 a_9698_2192.t6 VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X366 VSS.t151 saff_delay_unit_4/saff_2_0.nq a_10086_296# VSS.t150 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X367 saff_delay_unit_4/delay_unit_2_0.in_1.t0 saff_delay_unit_3/delay_unit_2_0.in_2.t17 VSS.t399 VSS.t398 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X368 saff_delay_unit_1/delay_unit_2_0.in_2.t2 start_pos.t8 VSS.t312 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X369 VDD.t5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 saff_delay_unit_0/saff_2_0.nq VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X370 a_14350_2192# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X371 a_9698_2192.t0 saff_delay_unit_5/delay_unit_2_0.in_1.t18 a_9786_2192# VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X372 a_10502_1376# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VDD.t172 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X373 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VDD.t315 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X374 VSS.t138 stop_strong.t47 a_7416_2192.t5 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X375 VSS.t15 a_15066_1376# saff_delay_unit_6/saff_2_0.nq VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X376 a_958_730# a_690_160# term_0.t2 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X377 VDD.t73 saff_delay_unit_7/delay_unit_2_0.in_1.t16 saff_delay_unit_7/delay_unit_2_0.in_2.t2 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X378 saff_delay_unit_6/delay_unit_2_0.in_1.t5 saff_delay_unit_5/delay_unit_2_0.in_2.t18 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X379 a_3656_1376# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VSS.t258 VSS.t257 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X380 VSS.t383 stop_strong.t48 a_570_2192.t4 VSS.t382 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X381 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 stop_strong.t49 VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X382 saff_delay_unit_4/saff_2_0.nq a_10502_1376# a_10464_730# VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X383 a_14262_2192.t0 saff_delay_unit_7/delay_unit_2_0.in_1.t17 a_14350_2192# VSS.t203 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X384 saff_delay_unit_2/delay_unit_2_0.in_2.t1 saff_delay_unit_1/delay_unit_2_0.in_1.t17 VSS.t108 VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X385 VDD.t273 saff_delay_unit_3/delay_unit_2_0.in_2.t18 saff_delay_unit_4/delay_unit_2_0.in_1.t3 VDD.t272 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X386 VDD.t238 start_pos.t9 saff_delay_unit_1/delay_unit_2_0.in_2.t5 VDD.t237 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X387 VDD.t218 saff_delay_unit_6/saff_2_0.nq a_14650_730# VDD.t217 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X388 a_5398_2192.t0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X389 saff_delay_unit_3/delay_unit_2_0.in_2.t3 saff_delay_unit_2/delay_unit_2_0.in_1.t19 VDD.t191 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X390 a_570_2192.t0 saff_delay_unit_1/delay_unit_2_0.in_1.t18 a_658_2192# VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X391 saff_delay_unit_5/delay_unit_2_0.in_1.t1 saff_delay_unit_4/delay_unit_2_0.in_2.t19 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X392 a_658_2192# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X393 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X394 VDD.t223 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 a_7536_160# VDD.t222 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X395 a_1336_730# term_0.t5 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X396 saff_delay_unit_7/saff_2_0.nd.t4 saff_delay_unit_7/delay_unit_2_0.in_1.t18 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X397 VDD.t127 saff_delay_unit_4/saff_2_0.nq a_10086_730# VDD.t126 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X398 a_7504_2192# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VSS.t298 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X399 a_15028_296# term_6.t4 VSS.t170 VSS.t169 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X400 a_16544_2192.t3 saff_delay_unit_7/saff_2_0.nd.t17 a_16808_2192.t3 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X401 VSS.t164 saff_delay_unit_3/delay_unit_2_0.in_1.t17 saff_delay_unit_4/delay_unit_2_0.in_2.t1 VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X402 VSS.t33 stop_strong.t50 a_14262_2192.t8 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X403 term_4.t0 a_9818_160# VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X404 VDD.t37 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X405 a_11980_2192.t6 stop_strong.t51 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X406 VDD.t269 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_6/saff_2_0.nq VDD.t268 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X407 a_5222_2192# saff_delay_unit_3/delay_unit_2_0.in_1.t18 a_5134_2192.t10 VSS.t165 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X408 VDD.t246 saff_delay_unit_1/delay_unit_2_0.in_2.t19 saff_delay_unit_2/delay_unit_2_0.in_1.t3 VDD.t245 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X409 a_3656_1376# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X410 VDD.t134 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X411 VDD.t264 saff_delay_unit_4/delay_unit_2_0.in_1.t18 saff_delay_unit_4/delay_unit_2_0.in_2.t7 VDD.t263 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X412 a_5222_2192# saff_delay_unit_3/delay_unit_2_0.in_1.t19 a_5134_2192.t9 VSS.t167 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X413 a_17348_1376# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VSS.t263 VSS.t262 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X414 delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.d.t19 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X415 a_16808_2192.t0 saff_delay_unit_7/saff_2_0.nd.t18 a_16544_2192.t0 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X416 saff_delay_unit_6/delay_unit_2_0.in_2.t4 saff_delay_unit_5/delay_unit_2_0.in_1.t19 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X417 VDD.t142 saff_delay_unit_4/delay_unit_2_0.in_1.t19 saff_delay_unit_5/delay_unit_2_0.in_2.t3 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X418 VSS.t50 stop_strong.t52 a_9698_2192.t5 VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X419 a_2940_2192# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X420 VSS.t147 saff_delay_unit_6/delay_unit_2_0.in_1.t19 saff_delay_unit_6/delay_unit_2_0.in_2.t0 VSS.t146 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X421 saff_delay_unit_1/delay_unit_2_0.in_1.t0 start_neg.t8 VSS.t172 VSS.t171 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X422 VSS.t297 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 a_14382_160# VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X423 VSS.t52 stop_strong.t53 a_9698_2192.t4 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X424 a_15028_730# term_6.t5 VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X425 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 a_12068_2192# VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X426 delay_unit_2_0.out_1.t3 saff_delay_unit_7/saff_2_0.nd.t19 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X427 VDD.t291 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X428 VSS.t212 a_8220_1376# saff_delay_unit_3/saff_2_0.nq VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X429 VDD.t67 start_neg.t9 start_pos.t0 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X430 term_4.t2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VDD.t287 VDD.t286 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X431 a_14526_2192.t0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VSS.t128 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X432 VSS.t327 stop_strong.t54 a_7416_2192.t4 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X433 saff_delay_unit_2/delay_unit_2_0.in_2.t0 saff_delay_unit_1/delay_unit_2_0.in_1.t19 VSS.t105 VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X434 VDD.t83 saff_delay_unit_3/delay_unit_2_0.in_2.t19 saff_delay_unit_3/delay_unit_2_0.in_1.t7 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X435 VSS.t335 saff_delay_unit_7/saff_2_0.nq a_16932_296# VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X436 VDD.t170 saff_delay_unit_7/delay_unit_2_0.in_1.t19 saff_delay_unit_7/saff_2_0.nd.t3 VDD.t169 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X437 a_12244_2192.t2 saff_delay_unit_6/delay_unit_2_0.in_2.t19 a_11980_2192.t12 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X438 VDD.t262 stop_strong.t55 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 VDD.t261 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X439 saff_delay_unit_6/delay_unit_2_0.in_1.t2 saff_delay_unit_5/delay_unit_2_0.in_2.t19 VSS.t200 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
R0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 890.727
R1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 742.783
R2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 665.16
R3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 623.388
R4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 523.774
R5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 431.807
R6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 427.875
R7 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 364.733
R8 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 208.5
R9 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 168.007
R10 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R11 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 31.2728
R12 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R13 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R14 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R15 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R16 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 8.00471
R17 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R18 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R19 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R20 VDD.n388 VDD.n72 2143.14
R21 VDD.n402 VDD.n64 2143.14
R22 VDD.n416 VDD.n56 2143.14
R23 VDD.n430 VDD.n48 2143.14
R24 VDD.n444 VDD.n40 2143.14
R25 VDD.n458 VDD.n32 2143.14
R26 VDD.n472 VDD.n24 2143.14
R27 VDD.n13 VDD.n7 2143.14
R28 VDD.n392 VDD.n387 2138.43
R29 VDD.n406 VDD.n401 2138.43
R30 VDD.n420 VDD.n415 2138.43
R31 VDD.n434 VDD.n429 2138.43
R32 VDD.n448 VDD.n443 2138.43
R33 VDD.n462 VDD.n457 2138.43
R34 VDD.n476 VDD.n471 2138.43
R35 VDD.n9 VDD.n8 2138.43
R36 VDD.n375 VDD.n373 2130.42
R37 VDD.n359 VDD.n357 2130.42
R38 VDD.n343 VDD.n341 2130.42
R39 VDD.n327 VDD.n325 2130.42
R40 VDD.n311 VDD.n309 2130.42
R41 VDD.n295 VDD.n293 2130.42
R42 VDD.n279 VDD.n277 2130.42
R43 VDD.n263 VDD.n261 2130.42
R44 VDD.n247 VDD.n245 2130.42
R45 VDD.n378 VDD.n374 2125.42
R46 VDD.n362 VDD.n358 2125.42
R47 VDD.n346 VDD.n342 2125.42
R48 VDD.n330 VDD.n326 2125.42
R49 VDD.n314 VDD.n310 2125.42
R50 VDD.n298 VDD.n294 2125.42
R51 VDD.n282 VDD.n278 2125.42
R52 VDD.n266 VDD.n262 2125.42
R53 VDD.n250 VDD.n246 2125.42
R54 VDD.n181 VDD.n179 1656.75
R55 VDD.n171 VDD.n169 1656.75
R56 VDD.n161 VDD.n159 1656.75
R57 VDD.n151 VDD.n149 1656.75
R58 VDD.n141 VDD.n139 1656.75
R59 VDD.n131 VDD.n129 1656.75
R60 VDD.n121 VDD.n119 1656.75
R61 VDD.n112 VDD.n110 1656.75
R62 VDD.n179 VDD.n178 1600.08
R63 VDD.n169 VDD.n168 1600.08
R64 VDD.n159 VDD.n158 1600.08
R65 VDD.n149 VDD.n148 1600.08
R66 VDD.n139 VDD.n138 1600.08
R67 VDD.n129 VDD.n128 1600.08
R68 VDD.n119 VDD.n118 1600.08
R69 VDD.n110 VDD.n109 1600.08
R70 VDD.n390 VDD.n387 1486.67
R71 VDD.n404 VDD.n401 1486.67
R72 VDD.n418 VDD.n415 1486.67
R73 VDD.n432 VDD.n429 1486.67
R74 VDD.n446 VDD.n443 1486.67
R75 VDD.n460 VDD.n457 1486.67
R76 VDD.n474 VDD.n471 1486.67
R77 VDD.n10 VDD.n8 1486.67
R78 VDD.n373 VDD.n193 1361.05
R79 VDD.n357 VDD.n199 1361.05
R80 VDD.n341 VDD.n205 1361.05
R81 VDD.n325 VDD.n211 1361.05
R82 VDD.n309 VDD.n217 1361.05
R83 VDD.n293 VDD.n223 1361.05
R84 VDD.n277 VDD.n229 1361.05
R85 VDD.n261 VDD.n235 1361.05
R86 VDD.n245 VDD.n241 1361.05
R87 VDD.n395 VDD.n69 228.601
R88 VDD.n409 VDD.n61 228.601
R89 VDD.n423 VDD.n53 228.601
R90 VDD.n437 VDD.n45 228.601
R91 VDD.n451 VDD.n37 228.601
R92 VDD.n465 VDD.n29 228.601
R93 VDD.n479 VDD.n21 228.601
R94 VDD.n15 VDD.n6 228.601
R95 VDD.n394 VDD.n393 228.1
R96 VDD.n408 VDD.n407 228.1
R97 VDD.n422 VDD.n421 228.1
R98 VDD.n436 VDD.n435 228.1
R99 VDD.n450 VDD.n449 228.1
R100 VDD.n464 VDD.n463 228.1
R101 VDD.n478 VDD.n477 228.1
R102 VDD.n14 VDD.n0 228.1
R103 VDD.n380 VDD.n372 227.244
R104 VDD.n364 VDD.n356 227.244
R105 VDD.n348 VDD.n340 227.244
R106 VDD.n332 VDD.n324 227.244
R107 VDD.n316 VDD.n308 227.244
R108 VDD.n300 VDD.n292 227.244
R109 VDD.n284 VDD.n276 227.244
R110 VDD.n268 VDD.n260 227.244
R111 VDD.n252 VDD.n244 227.244
R112 VDD.n379 VDD.n188 226.712
R113 VDD.n363 VDD.n194 226.712
R114 VDD.n347 VDD.n200 226.712
R115 VDD.n331 VDD.n206 226.712
R116 VDD.n315 VDD.n212 226.712
R117 VDD.n299 VDD.n218 226.712
R118 VDD.n283 VDD.n224 226.712
R119 VDD.n267 VDD.n230 226.712
R120 VDD.n251 VDD.n236 226.712
R121 VDD.n182 VDD.t36 196.429
R122 VDD.n172 VDD.t290 196.429
R123 VDD.n162 VDD.t209 196.429
R124 VDD.n152 VDD.t133 196.429
R125 VDD.n142 VDD.t302 196.429
R126 VDD.n132 VDD.t42 196.429
R127 VDD.n122 VDD.t179 196.429
R128 VDD.n113 VDD.t231 196.429
R129 VDD.n184 VDD.n178 186.093
R130 VDD.n174 VDD.n168 186.093
R131 VDD.n164 VDD.n158 186.093
R132 VDD.n154 VDD.n148 186.093
R133 VDD.n144 VDD.n138 186.093
R134 VDD.n134 VDD.n128 186.093
R135 VDD.n124 VDD.n118 186.093
R136 VDD.n115 VDD.n109 186.093
R137 VDD.n180 VDD.t137 183.929
R138 VDD.n170 VDD.t122 183.929
R139 VDD.n160 VDD.t30 183.929
R140 VDD.n150 VDD.t314 183.929
R141 VDD.n140 VDD.t118 183.929
R142 VDD.n130 VDD.t147 183.929
R143 VDD.n120 VDD.t149 183.929
R144 VDD.n111 VDD.t193 183.929
R145 VDD.n184 VDD.n77 176.72
R146 VDD.n174 VDD.n81 176.72
R147 VDD.n164 VDD.n85 176.72
R148 VDD.n154 VDD.n89 176.72
R149 VDD.n144 VDD.n93 176.72
R150 VDD.n134 VDD.n97 176.72
R151 VDD.n124 VDD.n101 176.72
R152 VDD.n115 VDD.n105 176.72
R153 VDD.t60 VDD.n388 169.983
R154 VDD.t102 VDD.n402 169.983
R155 VDD.t58 VDD.n416 169.983
R156 VDD.t26 VDD.n430 169.983
R157 VDD.t171 VDD.n444 169.983
R158 VDD.t96 VDD.n458 169.983
R159 VDD.t276 VDD.n472 169.983
R160 VDD.t197 VDD.n7 169.983
R161 VDD.n392 VDD.t292 164.046
R162 VDD.n406 VDD.t62 164.046
R163 VDD.n420 VDD.t229 164.046
R164 VDD.n434 VDD.t222 164.046
R165 VDD.n448 VDD.t90 164.046
R166 VDD.n462 VDD.t40 164.046
R167 VDD.n476 VDD.t70 164.046
R168 VDD.t235 VDD.n9 164.046
R169 VDD.n380 VDD.n193 160.596
R170 VDD.n364 VDD.n199 160.596
R171 VDD.n348 VDD.n205 160.596
R172 VDD.n332 VDD.n211 160.596
R173 VDD.n316 VDD.n217 160.596
R174 VDD.n300 VDD.n223 160.596
R175 VDD.n284 VDD.n229 160.596
R176 VDD.n268 VDD.n235 160.596
R177 VDD.n252 VDD.n241 160.596
R178 VDD.n394 VDD.n73 158.578
R179 VDD.n408 VDD.n65 158.578
R180 VDD.n422 VDD.n57 158.578
R181 VDD.n436 VDD.n49 158.578
R182 VDD.n450 VDD.n41 158.578
R183 VDD.n464 VDD.n33 158.578
R184 VDD.n478 VDD.n25 158.578
R185 VDD.n14 VDD.n2 158.578
R186 VDD.t241 VDD.n375 150.466
R187 VDD.t66 VDD.n374 150.466
R188 VDD.t76 VDD.n359 150.466
R189 VDD.t249 VDD.n358 150.466
R190 VDD.t177 VDD.n343 150.466
R191 VDD.t14 VDD.n342 150.466
R192 VDD.t112 VDD.n327 150.466
R193 VDD.t82 VDD.n326 150.466
R194 VDD.t184 VDD.n311 150.466
R195 VDD.t64 VDD.n310 150.466
R196 VDD.t225 VDD.n295 150.466
R197 VDD.t312 VDD.n294 150.466
R198 VDD.t145 VDD.n279 150.466
R199 VDD.t28 VDD.n278 150.466
R200 VDD.t298 VDD.n263 150.466
R201 VDD.t114 VDD.n262 150.466
R202 VDD.t166 VDD.n247 150.466
R203 VDD.t88 VDD.n246 150.466
R204 VDD.t153 VDD.n181 146.282
R205 VDD.t106 VDD.n171 146.282
R206 VDD.t173 VDD.n161 146.282
R207 VDD.t155 VDD.n151 146.282
R208 VDD.t92 VDD.n141 146.282
R209 VDD.t308 VDD.n131 146.282
R210 VDD.t8 VDD.n121 146.282
R211 VDD.t124 VDD.n112 146.282
R212 VDD.t278 VDD.n178 144.881
R213 VDD.t108 VDD.n168 144.881
R214 VDD.t213 VDD.n158 144.881
R215 VDD.t22 VDD.n148 144.881
R216 VDD.t20 VDD.n138 144.881
R217 VDD.t310 VDD.n128 144.881
R218 VDD.t261 VDD.n118 144.881
R219 VDD.t151 VDD.n109 144.881
R220 VDD.t294 VDD.n391 143.49
R221 VDD.t215 VDD.n405 143.49
R222 VDD.t46 VDD.n419 143.49
R223 VDD.t266 VDD.n433 143.49
R224 VDD.t126 VDD.n447 143.49
R225 VDD.t162 VDD.n461 143.49
R226 VDD.t217 VDD.n475 143.49
R227 VDD.n11 VDD.t270 143.49
R228 VDD.n389 VDD.t300 141.511
R229 VDD.n403 VDD.t51 141.511
R230 VDD.n417 VDD.t6 141.511
R231 VDD.n431 VDD.t49 141.511
R232 VDD.n445 VDD.t211 141.511
R233 VDD.n459 VDD.t207 141.511
R234 VDD.n473 VDD.t143 141.511
R235 VDD.n12 VDD.t18 141.511
R236 VDD.n376 VDD.t239 135.981
R237 VDD.n360 VDD.t80 135.981
R238 VDD.n344 VDD.t86 135.981
R239 VDD.n328 VDD.t199 135.981
R240 VDD.n312 VDD.t263 135.981
R241 VDD.n296 VDD.t282 135.981
R242 VDD.n280 VDD.t306 135.981
R243 VDD.n264 VDD.t72 135.981
R244 VDD.n248 VDD.t129 135.981
R245 VDD.n377 VDD.t274 132.256
R246 VDD.n361 VDD.t247 132.256
R247 VDD.n345 VDD.t16 132.256
R248 VDD.n329 VDD.t316 132.256
R249 VDD.n313 VDD.t54 132.256
R250 VDD.n297 VDD.t110 132.256
R251 VDD.n281 VDD.t56 132.256
R252 VDD.n265 VDD.t304 132.256
R253 VDD.n249 VDD.t32 132.256
R254 VDD.t4 VDD.t60 87.0838
R255 VDD.t44 VDD.t4 87.0838
R256 VDD.t300 VDD.t44 87.0838
R257 VDD.t45 VDD.t294 87.0838
R258 VDD.t259 VDD.t45 87.0838
R259 VDD.t292 VDD.t259 87.0838
R260 VDD.t104 VDD.t102 87.0838
R261 VDD.t53 VDD.t104 87.0838
R262 VDD.t51 VDD.t53 87.0838
R263 VDD.t48 VDD.t215 87.0838
R264 VDD.t139 VDD.t48 87.0838
R265 VDD.t62 VDD.t139 87.0838
R266 VDD.t94 VDD.t58 87.0838
R267 VDD.t159 VDD.t94 87.0838
R268 VDD.t6 VDD.t159 87.0838
R269 VDD.t224 VDD.t46 87.0838
R270 VDD.t205 VDD.t224 87.0838
R271 VDD.t229 VDD.t205 87.0838
R272 VDD.t181 VDD.t26 87.0838
R273 VDD.t168 VDD.t181 87.0838
R274 VDD.t49 VDD.t168 87.0838
R275 VDD.t158 VDD.t266 87.0838
R276 VDD.t253 VDD.t158 87.0838
R277 VDD.t222 VDD.t253 87.0838
R278 VDD.t135 VDD.t171 87.0838
R279 VDD.t128 VDD.t135 87.0838
R280 VDD.t211 VDD.t128 87.0838
R281 VDD.t13 VDD.t126 87.0838
R282 VDD.t286 VDD.t13 87.0838
R283 VDD.t90 VDD.t286 87.0838
R284 VDD.t38 VDD.t96 87.0838
R285 VDD.t221 VDD.t38 87.0838
R286 VDD.t207 VDD.t221 87.0838
R287 VDD.t157 VDD.t162 87.0838
R288 VDD.t120 VDD.t157 87.0838
R289 VDD.t40 VDD.t120 87.0838
R290 VDD.t268 VDD.t276 87.0838
R291 VDD.t10 VDD.t268 87.0838
R292 VDD.t143 VDD.t10 87.0838
R293 VDD.t183 VDD.t217 87.0838
R294 VDD.t164 VDD.t183 87.0838
R295 VDD.t70 VDD.t164 87.0838
R296 VDD.t233 VDD.t197 87.0838
R297 VDD.t192 VDD.t233 87.0838
R298 VDD.t18 VDD.t192 87.0838
R299 VDD.t270 VDD.t265 87.0838
R300 VDD.t265 VDD.t195 87.0838
R301 VDD.t195 VDD.t235 87.0838
R302 VDD.n78 VDD.t279 85.2064
R303 VDD.n82 VDD.t109 85.2064
R304 VDD.n86 VDD.t214 85.2064
R305 VDD.n90 VDD.t23 85.2064
R306 VDD.n94 VDD.t21 85.2064
R307 VDD.n98 VDD.t311 85.2064
R308 VDD.n102 VDD.t262 85.2064
R309 VDD.n106 VDD.t152 85.2064
R310 VDD.n75 VDD.t295 85.0216
R311 VDD.n397 VDD.t301 85.0216
R312 VDD.n67 VDD.t216 85.0216
R313 VDD.n411 VDD.t52 85.0216
R314 VDD.n59 VDD.t47 85.0216
R315 VDD.n425 VDD.t7 85.0216
R316 VDD.n51 VDD.t267 85.0216
R317 VDD.n439 VDD.t50 85.0216
R318 VDD.n43 VDD.t127 85.0216
R319 VDD.n453 VDD.t212 85.0216
R320 VDD.n35 VDD.t163 85.0216
R321 VDD.n467 VDD.t208 85.0216
R322 VDD.n27 VDD.t218 85.0216
R323 VDD.n481 VDD.t144 85.0216
R324 VDD.n18 VDD.t271 85.0216
R325 VDD.n3 VDD.t19 85.0216
R326 VDD.n80 VDD.t154 84.7281
R327 VDD.n79 VDD.t37 84.7281
R328 VDD.n78 VDD.t138 84.7281
R329 VDD.n84 VDD.t107 84.7281
R330 VDD.n83 VDD.t291 84.7281
R331 VDD.n82 VDD.t123 84.7281
R332 VDD.n88 VDD.t174 84.7281
R333 VDD.n87 VDD.t210 84.7281
R334 VDD.n86 VDD.t31 84.7281
R335 VDD.n92 VDD.t156 84.7281
R336 VDD.n91 VDD.t134 84.7281
R337 VDD.n90 VDD.t315 84.7281
R338 VDD.n96 VDD.t93 84.7281
R339 VDD.n95 VDD.t303 84.7281
R340 VDD.n94 VDD.t119 84.7281
R341 VDD.n100 VDD.t309 84.7281
R342 VDD.n99 VDD.t43 84.7281
R343 VDD.n98 VDD.t148 84.7281
R344 VDD.n104 VDD.t9 84.7281
R345 VDD.n103 VDD.t180 84.7281
R346 VDD.n102 VDD.t150 84.7281
R347 VDD.n108 VDD.t125 84.7281
R348 VDD.n107 VDD.t232 84.7281
R349 VDD.n106 VDD.t194 84.7281
R350 VDD.t237 VDD.t241 81.9613
R351 VDD.t243 VDD.t237 81.9613
R352 VDD.t239 VDD.t243 81.9613
R353 VDD.t274 VDD.t201 81.9613
R354 VDD.t201 VDD.t280 81.9613
R355 VDD.t280 VDD.t66 81.9613
R356 VDD.t78 VDD.t76 81.9613
R357 VDD.t74 VDD.t78 81.9613
R358 VDD.t80 VDD.t74 81.9613
R359 VDD.t247 VDD.t245 81.9613
R360 VDD.t245 VDD.t251 81.9613
R361 VDD.t251 VDD.t249 81.9613
R362 VDD.t84 VDD.t177 81.9613
R363 VDD.t190 VDD.t84 81.9613
R364 VDD.t86 VDD.t190 81.9613
R365 VDD.t16 VDD.t0 81.9613
R366 VDD.t0 VDD.t2 81.9613
R367 VDD.t2 VDD.t14 81.9613
R368 VDD.t188 VDD.t112 81.9613
R369 VDD.t219 VDD.t188 81.9613
R370 VDD.t199 VDD.t219 81.9613
R371 VDD.t316 VDD.t272 81.9613
R372 VDD.t272 VDD.t318 81.9613
R373 VDD.t318 VDD.t82 81.9613
R374 VDD.t141 VDD.t184 81.9613
R375 VDD.t203 VDD.t141 81.9613
R376 VDD.t263 VDD.t203 81.9613
R377 VDD.t54 VDD.t24 81.9613
R378 VDD.t24 VDD.t175 81.9613
R379 VDD.t175 VDD.t64 81.9613
R380 VDD.t296 VDD.t225 81.9613
R381 VDD.t227 VDD.t296 81.9613
R382 VDD.t282 VDD.t227 81.9613
R383 VDD.t110 VDD.t131 81.9613
R384 VDD.t131 VDD.t284 81.9613
R385 VDD.t284 VDD.t312 81.9613
R386 VDD.t100 VDD.t145 81.9613
R387 VDD.t257 VDD.t100 81.9613
R388 VDD.t306 VDD.t257 81.9613
R389 VDD.t56 VDD.t98 81.9613
R390 VDD.t98 VDD.t160 81.9613
R391 VDD.t160 VDD.t28 81.9613
R392 VDD.t169 VDD.t298 81.9613
R393 VDD.t186 VDD.t169 81.9613
R394 VDD.t72 VDD.t186 81.9613
R395 VDD.t304 VDD.t288 81.9613
R396 VDD.t288 VDD.t34 81.9613
R397 VDD.t34 VDD.t114 81.9613
R398 VDD.t68 VDD.t166 81.9613
R399 VDD.t11 VDD.t68 81.9613
R400 VDD.t129 VDD.t11 81.9613
R401 VDD.t32 VDD.t255 81.9613
R402 VDD.t255 VDD.t116 81.9613
R403 VDD.t116 VDD.t88 81.9613
R404 VDD.t137 VDD.t278 78.5719
R405 VDD.t36 VDD.t153 78.5719
R406 VDD.t122 VDD.t108 78.5719
R407 VDD.t290 VDD.t106 78.5719
R408 VDD.t30 VDD.t213 78.5719
R409 VDD.t209 VDD.t173 78.5719
R410 VDD.t314 VDD.t22 78.5719
R411 VDD.t133 VDD.t155 78.5719
R412 VDD.t118 VDD.t20 78.5719
R413 VDD.t302 VDD.t92 78.5719
R414 VDD.t147 VDD.t310 78.5719
R415 VDD.t42 VDD.t308 78.5719
R416 VDD.t149 VDD.t261 78.5719
R417 VDD.t179 VDD.t8 78.5719
R418 VDD.t193 VDD.t151 78.5719
R419 VDD.t231 VDD.t124 78.5719
R420 VDD.n383 VDD.n189 75.7173
R421 VDD.n382 VDD.n190 75.7173
R422 VDD.n192 VDD.n191 75.7173
R423 VDD.n370 VDD.n369 75.7173
R424 VDD.n367 VDD.n195 75.7173
R425 VDD.n366 VDD.n196 75.7173
R426 VDD.n198 VDD.n197 75.7173
R427 VDD.n354 VDD.n353 75.7173
R428 VDD.n351 VDD.n201 75.7173
R429 VDD.n350 VDD.n202 75.7173
R430 VDD.n204 VDD.n203 75.7173
R431 VDD.n338 VDD.n337 75.7173
R432 VDD.n335 VDD.n207 75.7173
R433 VDD.n334 VDD.n208 75.7173
R434 VDD.n210 VDD.n209 75.7173
R435 VDD.n322 VDD.n321 75.7173
R436 VDD.n319 VDD.n213 75.7173
R437 VDD.n318 VDD.n214 75.7173
R438 VDD.n216 VDD.n215 75.7173
R439 VDD.n306 VDD.n305 75.7173
R440 VDD.n303 VDD.n219 75.7173
R441 VDD.n302 VDD.n220 75.7173
R442 VDD.n222 VDD.n221 75.7173
R443 VDD.n290 VDD.n289 75.7173
R444 VDD.n287 VDD.n225 75.7173
R445 VDD.n286 VDD.n226 75.7173
R446 VDD.n228 VDD.n227 75.7173
R447 VDD.n274 VDD.n273 75.7173
R448 VDD.n271 VDD.n231 75.7173
R449 VDD.n270 VDD.n232 75.7173
R450 VDD.n234 VDD.n233 75.7173
R451 VDD.n258 VDD.n257 75.7173
R452 VDD.n255 VDD.n237 75.7173
R453 VDD.n254 VDD.n238 75.7173
R454 VDD.n240 VDD.n239 75.7173
R455 VDD.n243 VDD.n242 75.7173
R456 VDD.n76 VDD.n74 75.5
R457 VDD.n398 VDD.n70 75.5
R458 VDD.n68 VDD.n66 75.5
R459 VDD.n412 VDD.n62 75.5
R460 VDD.n60 VDD.n58 75.5
R461 VDD.n426 VDD.n54 75.5
R462 VDD.n52 VDD.n50 75.5
R463 VDD.n440 VDD.n46 75.5
R464 VDD.n44 VDD.n42 75.5
R465 VDD.n454 VDD.n38 75.5
R466 VDD.n36 VDD.n34 75.5
R467 VDD.n468 VDD.n30 75.5
R468 VDD.n28 VDD.n26 75.5
R469 VDD.n482 VDD.n22 75.5
R470 VDD.n19 VDD.n1 75.5
R471 VDD.n5 VDD.n4 75.5
R472 VDD.n183 VDD.n182 38.0519
R473 VDD.n173 VDD.n172 38.0519
R474 VDD.n163 VDD.n162 38.0519
R475 VDD.n153 VDD.n152 38.0519
R476 VDD.n143 VDD.n142 38.0519
R477 VDD.n133 VDD.n132 38.0519
R478 VDD.n123 VDD.n122 38.0519
R479 VDD.n114 VDD.n113 38.0519
R480 VDD.n393 VDD.n392 20.5561
R481 VDD.n390 VDD.n73 20.5561
R482 VDD.n391 VDD.n390 20.5561
R483 VDD.n388 VDD.n69 20.5561
R484 VDD.n407 VDD.n406 20.5561
R485 VDD.n404 VDD.n65 20.5561
R486 VDD.n405 VDD.n404 20.5561
R487 VDD.n402 VDD.n61 20.5561
R488 VDD.n421 VDD.n420 20.5561
R489 VDD.n418 VDD.n57 20.5561
R490 VDD.n419 VDD.n418 20.5561
R491 VDD.n416 VDD.n53 20.5561
R492 VDD.n435 VDD.n434 20.5561
R493 VDD.n432 VDD.n49 20.5561
R494 VDD.n433 VDD.n432 20.5561
R495 VDD.n430 VDD.n45 20.5561
R496 VDD.n449 VDD.n448 20.5561
R497 VDD.n446 VDD.n41 20.5561
R498 VDD.n447 VDD.n446 20.5561
R499 VDD.n444 VDD.n37 20.5561
R500 VDD.n463 VDD.n462 20.5561
R501 VDD.n460 VDD.n33 20.5561
R502 VDD.n461 VDD.n460 20.5561
R503 VDD.n458 VDD.n29 20.5561
R504 VDD.n477 VDD.n476 20.5561
R505 VDD.n474 VDD.n25 20.5561
R506 VDD.n475 VDD.n474 20.5561
R507 VDD.n472 VDD.n21 20.5561
R508 VDD.n9 VDD.n0 20.5561
R509 VDD.n10 VDD.n2 20.5561
R510 VDD.n11 VDD.n10 20.5561
R511 VDD.n7 VDD.n6 20.5561
R512 VDD.n181 VDD.n77 16.8187
R513 VDD.n171 VDD.n81 16.8187
R514 VDD.n161 VDD.n85 16.8187
R515 VDD.n151 VDD.n89 16.8187
R516 VDD.n141 VDD.n93 16.8187
R517 VDD.n131 VDD.n97 16.8187
R518 VDD.n121 VDD.n101 16.8187
R519 VDD.n112 VDD.n105 16.8187
R520 VDD.n376 VDD.n193 15.4172
R521 VDD.n374 VDD.n188 15.4172
R522 VDD.n375 VDD.n372 15.4172
R523 VDD.n360 VDD.n199 15.4172
R524 VDD.n358 VDD.n194 15.4172
R525 VDD.n359 VDD.n356 15.4172
R526 VDD.n344 VDD.n205 15.4172
R527 VDD.n342 VDD.n200 15.4172
R528 VDD.n343 VDD.n340 15.4172
R529 VDD.n328 VDD.n211 15.4172
R530 VDD.n326 VDD.n206 15.4172
R531 VDD.n327 VDD.n324 15.4172
R532 VDD.n312 VDD.n217 15.4172
R533 VDD.n310 VDD.n212 15.4172
R534 VDD.n311 VDD.n308 15.4172
R535 VDD.n296 VDD.n223 15.4172
R536 VDD.n294 VDD.n218 15.4172
R537 VDD.n295 VDD.n292 15.4172
R538 VDD.n280 VDD.n229 15.4172
R539 VDD.n278 VDD.n224 15.4172
R540 VDD.n279 VDD.n276 15.4172
R541 VDD.n264 VDD.n235 15.4172
R542 VDD.n262 VDD.n230 15.4172
R543 VDD.n263 VDD.n260 15.4172
R544 VDD.n248 VDD.n241 15.4172
R545 VDD.n246 VDD.n236 15.4172
R546 VDD.n247 VDD.n244 15.4172
R547 VDD.n182 VDD.n180 12.5005
R548 VDD.n172 VDD.n170 12.5005
R549 VDD.n162 VDD.n160 12.5005
R550 VDD.n152 VDD.n150 12.5005
R551 VDD.n142 VDD.n140 12.5005
R552 VDD.n132 VDD.n130 12.5005
R553 VDD.n122 VDD.n120 12.5005
R554 VDD.n113 VDD.n111 12.5005
R555 VDD.n379 VDD.n378 11.563
R556 VDD.n378 VDD.n377 11.563
R557 VDD.n363 VDD.n362 11.563
R558 VDD.n362 VDD.n361 11.563
R559 VDD.n347 VDD.n346 11.563
R560 VDD.n346 VDD.n345 11.563
R561 VDD.n331 VDD.n330 11.563
R562 VDD.n330 VDD.n329 11.563
R563 VDD.n315 VDD.n314 11.563
R564 VDD.n314 VDD.n313 11.563
R565 VDD.n299 VDD.n298 11.563
R566 VDD.n298 VDD.n297 11.563
R567 VDD.n283 VDD.n282 11.563
R568 VDD.n282 VDD.n281 11.563
R569 VDD.n267 VDD.n266 11.563
R570 VDD.n266 VDD.n265 11.563
R571 VDD.n251 VDD.n250 11.563
R572 VDD.n250 VDD.n249 11.563
R573 VDD.n189 VDD.t281 9.52217
R574 VDD.n189 VDD.t67 9.52217
R575 VDD.n190 VDD.t275 9.52217
R576 VDD.n190 VDD.t202 9.52217
R577 VDD.n191 VDD.t244 9.52217
R578 VDD.n191 VDD.t240 9.52217
R579 VDD.n369 VDD.t242 9.52217
R580 VDD.n369 VDD.t238 9.52217
R581 VDD.n195 VDD.t252 9.52217
R582 VDD.n195 VDD.t250 9.52217
R583 VDD.n196 VDD.t248 9.52217
R584 VDD.n196 VDD.t246 9.52217
R585 VDD.n197 VDD.t75 9.52217
R586 VDD.n197 VDD.t81 9.52217
R587 VDD.n353 VDD.t77 9.52217
R588 VDD.n353 VDD.t79 9.52217
R589 VDD.n201 VDD.t3 9.52217
R590 VDD.n201 VDD.t15 9.52217
R591 VDD.n202 VDD.t17 9.52217
R592 VDD.n202 VDD.t1 9.52217
R593 VDD.n203 VDD.t191 9.52217
R594 VDD.n203 VDD.t87 9.52217
R595 VDD.n337 VDD.t178 9.52217
R596 VDD.n337 VDD.t85 9.52217
R597 VDD.n207 VDD.t319 9.52217
R598 VDD.n207 VDD.t83 9.52217
R599 VDD.n208 VDD.t317 9.52217
R600 VDD.n208 VDD.t273 9.52217
R601 VDD.n209 VDD.t220 9.52217
R602 VDD.n209 VDD.t200 9.52217
R603 VDD.n321 VDD.t113 9.52217
R604 VDD.n321 VDD.t189 9.52217
R605 VDD.n213 VDD.t176 9.52217
R606 VDD.n213 VDD.t65 9.52217
R607 VDD.n214 VDD.t55 9.52217
R608 VDD.n214 VDD.t25 9.52217
R609 VDD.n215 VDD.t204 9.52217
R610 VDD.n215 VDD.t264 9.52217
R611 VDD.n305 VDD.t185 9.52217
R612 VDD.n305 VDD.t142 9.52217
R613 VDD.n219 VDD.t285 9.52217
R614 VDD.n219 VDD.t313 9.52217
R615 VDD.n220 VDD.t111 9.52217
R616 VDD.n220 VDD.t132 9.52217
R617 VDD.n221 VDD.t228 9.52217
R618 VDD.n221 VDD.t283 9.52217
R619 VDD.n289 VDD.t226 9.52217
R620 VDD.n289 VDD.t297 9.52217
R621 VDD.n225 VDD.t161 9.52217
R622 VDD.n225 VDD.t29 9.52217
R623 VDD.n226 VDD.t57 9.52217
R624 VDD.n226 VDD.t99 9.52217
R625 VDD.n227 VDD.t258 9.52217
R626 VDD.n227 VDD.t307 9.52217
R627 VDD.n273 VDD.t146 9.52217
R628 VDD.n273 VDD.t101 9.52217
R629 VDD.n231 VDD.t35 9.52217
R630 VDD.n231 VDD.t115 9.52217
R631 VDD.n232 VDD.t305 9.52217
R632 VDD.n232 VDD.t289 9.52217
R633 VDD.n233 VDD.t187 9.52217
R634 VDD.n233 VDD.t73 9.52217
R635 VDD.n257 VDD.t299 9.52217
R636 VDD.n257 VDD.t170 9.52217
R637 VDD.n237 VDD.t117 9.52217
R638 VDD.n237 VDD.t89 9.52217
R639 VDD.n238 VDD.t33 9.52217
R640 VDD.n238 VDD.t256 9.52217
R641 VDD.n239 VDD.t12 9.52217
R642 VDD.n239 VDD.t130 9.52217
R643 VDD.n242 VDD.t167 9.52217
R644 VDD.n242 VDD.t69 9.52217
R645 VDD.n74 VDD.t260 9.52217
R646 VDD.n74 VDD.t293 9.52217
R647 VDD.n70 VDD.t61 9.52217
R648 VDD.n70 VDD.t5 9.52217
R649 VDD.n66 VDD.t140 9.52217
R650 VDD.n66 VDD.t63 9.52217
R651 VDD.n62 VDD.t103 9.52217
R652 VDD.n62 VDD.t105 9.52217
R653 VDD.n58 VDD.t206 9.52217
R654 VDD.n58 VDD.t230 9.52217
R655 VDD.n54 VDD.t59 9.52217
R656 VDD.n54 VDD.t95 9.52217
R657 VDD.n50 VDD.t254 9.52217
R658 VDD.n50 VDD.t223 9.52217
R659 VDD.n46 VDD.t27 9.52217
R660 VDD.n46 VDD.t182 9.52217
R661 VDD.n42 VDD.t287 9.52217
R662 VDD.n42 VDD.t91 9.52217
R663 VDD.n38 VDD.t172 9.52217
R664 VDD.n38 VDD.t136 9.52217
R665 VDD.n34 VDD.t121 9.52217
R666 VDD.n34 VDD.t41 9.52217
R667 VDD.n30 VDD.t97 9.52217
R668 VDD.n30 VDD.t39 9.52217
R669 VDD.n26 VDD.t165 9.52217
R670 VDD.n26 VDD.t71 9.52217
R671 VDD.n22 VDD.t277 9.52217
R672 VDD.n22 VDD.t269 9.52217
R673 VDD.n1 VDD.t196 9.52217
R674 VDD.n1 VDD.t236 9.52217
R675 VDD.n4 VDD.t198 9.52217
R676 VDD.n4 VDD.t234 9.52217
R677 VDD.n180 VDD.n179 6.60764
R678 VDD.n170 VDD.n169 6.60764
R679 VDD.n160 VDD.n159 6.60764
R680 VDD.n150 VDD.n149 6.60764
R681 VDD.n140 VDD.n139 6.60764
R682 VDD.n130 VDD.n129 6.60764
R683 VDD.n120 VDD.n119 6.60764
R684 VDD.n111 VDD.n110 6.60764
R685 VDD.n183 VDD.n179 5.77063
R686 VDD.n173 VDD.n169 5.77063
R687 VDD.n163 VDD.n159 5.77063
R688 VDD.n153 VDD.n149 5.77063
R689 VDD.n143 VDD.n139 5.77063
R690 VDD.n133 VDD.n129 5.77063
R691 VDD.n123 VDD.n119 5.77063
R692 VDD.n114 VDD.n110 5.77063
R693 VDD.n395 VDD.n72 5.44168
R694 VDD.n389 VDD.n72 5.44168
R695 VDD.n409 VDD.n64 5.44168
R696 VDD.n403 VDD.n64 5.44168
R697 VDD.n423 VDD.n56 5.44168
R698 VDD.n417 VDD.n56 5.44168
R699 VDD.n437 VDD.n48 5.44168
R700 VDD.n431 VDD.n48 5.44168
R701 VDD.n451 VDD.n40 5.44168
R702 VDD.n445 VDD.n40 5.44168
R703 VDD.n465 VDD.n32 5.44168
R704 VDD.n459 VDD.n32 5.44168
R705 VDD.n479 VDD.n24 5.44168
R706 VDD.n473 VDD.n24 5.44168
R707 VDD.n15 VDD.n13 5.44168
R708 VDD.n13 VDD.n12 5.44168
R709 VDD.n378 VDD.n373 5.0005
R710 VDD.n362 VDD.n357 5.0005
R711 VDD.n346 VDD.n341 5.0005
R712 VDD.n330 VDD.n325 5.0005
R713 VDD.n314 VDD.n309 5.0005
R714 VDD.n298 VDD.n293 5.0005
R715 VDD.n282 VDD.n277 5.0005
R716 VDD.n266 VDD.n261 5.0005
R717 VDD.n250 VDD.n245 5.0005
R718 VDD.n377 VDD.n376 3.72599
R719 VDD.n361 VDD.n360 3.72599
R720 VDD.n345 VDD.n344 3.72599
R721 VDD.n329 VDD.n328 3.72599
R722 VDD.n313 VDD.n312 3.72599
R723 VDD.n297 VDD.n296 3.72599
R724 VDD.n281 VDD.n280 3.72599
R725 VDD.n265 VDD.n264 3.72599
R726 VDD.n249 VDD.n248 3.72599
R727 VDD VDD.n385 3.03187
R728 VDD.n6 VDD.n5 2.56343
R729 VDD.n387 VDD.n72 2.35344
R730 VDD.n401 VDD.n64 2.35344
R731 VDD.n415 VDD.n56 2.35344
R732 VDD.n429 VDD.n48 2.35344
R733 VDD.n443 VDD.n40 2.35344
R734 VDD.n457 VDD.n32 2.35344
R735 VDD.n471 VDD.n24 2.35344
R736 VDD.n13 VDD.n8 2.35344
R737 VDD.n393 VDD.n386 2.32446
R738 VDD.n73 VDD.n71 2.32446
R739 VDD.n399 VDD.n69 2.32446
R740 VDD.n407 VDD.n400 2.32446
R741 VDD.n65 VDD.n63 2.32446
R742 VDD.n413 VDD.n61 2.32446
R743 VDD.n421 VDD.n414 2.32446
R744 VDD.n57 VDD.n55 2.32446
R745 VDD.n427 VDD.n53 2.32446
R746 VDD.n435 VDD.n428 2.32446
R747 VDD.n49 VDD.n47 2.32446
R748 VDD.n441 VDD.n45 2.32446
R749 VDD.n449 VDD.n442 2.32446
R750 VDD.n41 VDD.n39 2.32446
R751 VDD.n455 VDD.n37 2.32446
R752 VDD.n463 VDD.n456 2.32446
R753 VDD.n33 VDD.n31 2.32446
R754 VDD.n469 VDD.n29 2.32446
R755 VDD.n477 VDD.n470 2.32446
R756 VDD.n25 VDD.n23 2.32446
R757 VDD.n483 VDD.n21 2.32446
R758 VDD.n20 VDD.n0 2.32446
R759 VDD.n17 VDD.n2 2.32446
R760 VDD.n244 VDD.n243 2.21444
R761 VDD.n391 VDD.n389 1.97967
R762 VDD.n405 VDD.n403 1.97967
R763 VDD.n419 VDD.n417 1.97967
R764 VDD.n433 VDD.n431 1.97967
R765 VDD.n447 VDD.n445 1.97967
R766 VDD.n461 VDD.n459 1.97967
R767 VDD.n475 VDD.n473 1.97967
R768 VDD.n12 VDD.n11 1.97967
R769 VDD.n384 VDD.n188 1.96835
R770 VDD.n372 VDD.n371 1.96835
R771 VDD.n368 VDD.n194 1.96835
R772 VDD.n356 VDD.n355 1.96835
R773 VDD.n352 VDD.n200 1.96835
R774 VDD.n340 VDD.n339 1.96835
R775 VDD.n336 VDD.n206 1.96835
R776 VDD.n324 VDD.n323 1.96835
R777 VDD.n320 VDD.n212 1.96835
R778 VDD.n308 VDD.n307 1.96835
R779 VDD.n304 VDD.n218 1.96835
R780 VDD.n292 VDD.n291 1.96835
R781 VDD.n288 VDD.n224 1.96835
R782 VDD.n276 VDD.n275 1.96835
R783 VDD.n272 VDD.n230 1.96835
R784 VDD.n260 VDD.n259 1.96835
R785 VDD.n256 VDD.n236 1.96835
R786 VDD.n187 VDD.n77 1.92668
R787 VDD.n177 VDD.n81 1.92668
R788 VDD.n167 VDD.n85 1.92668
R789 VDD.n157 VDD.n89 1.92668
R790 VDD.n147 VDD.n93 1.92668
R791 VDD.n137 VDD.n97 1.92668
R792 VDD.n127 VDD.n101 1.92668
R793 VDD.n117 VDD.n105 1.92668
R794 VDD.n259 VDD 1.45623
R795 VDD.n275 VDD 1.45623
R796 VDD.n291 VDD 1.45623
R797 VDD.n307 VDD 1.45623
R798 VDD.n323 VDD 1.45623
R799 VDD.n339 VDD 1.45623
R800 VDD.n355 VDD 1.45623
R801 VDD.n371 VDD 1.45623
R802 VDD.n385 VDD 1.42472
R803 VDD.n125 VDD 1.04243
R804 VDD.n135 VDD 1.04243
R805 VDD.n145 VDD 1.04243
R806 VDD.n155 VDD 1.04243
R807 VDD.n165 VDD 1.04243
R808 VDD.n175 VDD 1.04243
R809 VDD.n185 VDD 1.04243
R810 VDD.n79 VDD.n78 0.957022
R811 VDD.n83 VDD.n82 0.957022
R812 VDD.n87 VDD.n86 0.957022
R813 VDD.n91 VDD.n90 0.957022
R814 VDD.n95 VDD.n94 0.957022
R815 VDD.n99 VDD.n98 0.957022
R816 VDD.n103 VDD.n102 0.957022
R817 VDD.n107 VDD.n106 0.957022
R818 VDD.n184 VDD.n183 0.713588
R819 VDD.n174 VDD.n173 0.713588
R820 VDD.n164 VDD.n163 0.713588
R821 VDD.n154 VDD.n153 0.713588
R822 VDD.n144 VDD.n143 0.713588
R823 VDD.n134 VDD.n133 0.713588
R824 VDD.n124 VDD.n123 0.713588
R825 VDD.n115 VDD.n114 0.713588
R826 VDD VDD.n483 0.669618
R827 VDD VDD.n469 0.669618
R828 VDD VDD.n455 0.669618
R829 VDD VDD.n441 0.669618
R830 VDD VDD.n427 0.669618
R831 VDD VDD.n413 0.669618
R832 VDD VDD.n399 0.669618
R833 VDD.n116 VDD.n115 0.647749
R834 VDD.n253 VDD.n252 0.58175
R835 VDD.n269 VDD.n268 0.58175
R836 VDD.n285 VDD.n284 0.58175
R837 VDD.n301 VDD.n300 0.58175
R838 VDD.n317 VDD.n316 0.58175
R839 VDD.n333 VDD.n332 0.58175
R840 VDD.n349 VDD.n348 0.58175
R841 VDD.n365 VDD.n364 0.58175
R842 VDD.n381 VDD.n380 0.58175
R843 VDD.n16 VDD.n15 0.58175
R844 VDD.n480 VDD.n479 0.58175
R845 VDD.n466 VDD.n465 0.58175
R846 VDD.n452 VDD.n451 0.58175
R847 VDD.n438 VDD.n437 0.58175
R848 VDD.n424 VDD.n423 0.58175
R849 VDD.n410 VDD.n409 0.58175
R850 VDD.n396 VDD.n395 0.58175
R851 VDD.n380 VDD.n379 0.533833
R852 VDD.n364 VDD.n363 0.533833
R853 VDD.n348 VDD.n347 0.533833
R854 VDD.n332 VDD.n331 0.533833
R855 VDD.n316 VDD.n315 0.533833
R856 VDD.n300 VDD.n299 0.533833
R857 VDD.n284 VDD.n283 0.533833
R858 VDD.n268 VDD.n267 0.533833
R859 VDD.n252 VDD.n251 0.533833
R860 VDD.n80 VDD.n79 0.478761
R861 VDD.n84 VDD.n83 0.478761
R862 VDD.n88 VDD.n87 0.478761
R863 VDD.n92 VDD.n91 0.478761
R864 VDD.n96 VDD.n95 0.478761
R865 VDD.n100 VDD.n99 0.478761
R866 VDD.n104 VDD.n103 0.478761
R867 VDD.n108 VDD.n107 0.478761
R868 VDD VDD.n117 0.394487
R869 VDD VDD.n127 0.394487
R870 VDD VDD.n137 0.394487
R871 VDD VDD.n147 0.394487
R872 VDD VDD.n157 0.394487
R873 VDD VDD.n167 0.394487
R874 VDD VDD.n177 0.394487
R875 VDD VDD.n187 0.394487
R876 VDD.n125 VDD.n124 0.358192
R877 VDD.n135 VDD.n134 0.358192
R878 VDD.n145 VDD.n144 0.358192
R879 VDD.n155 VDD.n154 0.358192
R880 VDD.n165 VDD.n164 0.358192
R881 VDD.n175 VDD.n174 0.358192
R882 VDD.n185 VDD.n184 0.358192
R883 VDD.n186 VDD.n80 0.337457
R884 VDD.n176 VDD.n84 0.337457
R885 VDD.n166 VDD.n88 0.337457
R886 VDD.n156 VDD.n92 0.337457
R887 VDD.n146 VDD.n96 0.337457
R888 VDD.n136 VDD.n100 0.337457
R889 VDD.n126 VDD.n104 0.337457
R890 VDD.n116 VDD.n108 0.337457
R891 VDD.n5 VDD.n3 0.324029
R892 VDD.n19 VDD.n18 0.324029
R893 VDD.n482 VDD.n481 0.324029
R894 VDD.n28 VDD.n27 0.324029
R895 VDD.n468 VDD.n467 0.324029
R896 VDD.n36 VDD.n35 0.324029
R897 VDD.n454 VDD.n453 0.324029
R898 VDD.n44 VDD.n43 0.324029
R899 VDD.n440 VDD.n439 0.324029
R900 VDD.n52 VDD.n51 0.324029
R901 VDD.n426 VDD.n425 0.324029
R902 VDD.n60 VDD.n59 0.324029
R903 VDD.n412 VDD.n411 0.324029
R904 VDD.n68 VDD.n67 0.324029
R905 VDD.n398 VDD.n397 0.324029
R906 VDD.n76 VDD.n75 0.324029
R907 VDD.n126 VDD.n125 0.290057
R908 VDD.n136 VDD.n135 0.290057
R909 VDD.n146 VDD.n145 0.290057
R910 VDD.n156 VDD.n155 0.290057
R911 VDD.n166 VDD.n165 0.290057
R912 VDD.n176 VDD.n175 0.290057
R913 VDD.n186 VDD.n185 0.290057
R914 VDD.n385 VDD 0.278981
R915 VDD.n395 VDD.n394 0.25148
R916 VDD.n409 VDD.n408 0.25148
R917 VDD.n423 VDD.n422 0.25148
R918 VDD.n437 VDD.n436 0.25148
R919 VDD.n451 VDD.n450 0.25148
R920 VDD.n465 VDD.n464 0.25148
R921 VDD.n479 VDD.n478 0.25148
R922 VDD.n15 VDD.n14 0.25148
R923 VDD.n253 VDD.n240 0.247896
R924 VDD.n254 VDD.n253 0.247896
R925 VDD.n269 VDD.n234 0.247896
R926 VDD.n270 VDD.n269 0.247896
R927 VDD.n285 VDD.n228 0.247896
R928 VDD.n286 VDD.n285 0.247896
R929 VDD.n301 VDD.n222 0.247896
R930 VDD.n302 VDD.n301 0.247896
R931 VDD.n317 VDD.n216 0.247896
R932 VDD.n318 VDD.n317 0.247896
R933 VDD.n333 VDD.n210 0.247896
R934 VDD.n334 VDD.n333 0.247896
R935 VDD.n349 VDD.n204 0.247896
R936 VDD.n350 VDD.n349 0.247896
R937 VDD.n365 VDD.n198 0.247896
R938 VDD.n366 VDD.n365 0.247896
R939 VDD.n381 VDD.n192 0.247896
R940 VDD.n382 VDD.n381 0.247896
R941 VDD.n256 VDD.n255 0.246594
R942 VDD.n259 VDD.n258 0.246594
R943 VDD.n272 VDD.n271 0.246594
R944 VDD.n275 VDD.n274 0.246594
R945 VDD.n288 VDD.n287 0.246594
R946 VDD.n291 VDD.n290 0.246594
R947 VDD.n304 VDD.n303 0.246594
R948 VDD.n307 VDD.n306 0.246594
R949 VDD.n320 VDD.n319 0.246594
R950 VDD.n323 VDD.n322 0.246594
R951 VDD.n336 VDD.n335 0.246594
R952 VDD.n339 VDD.n338 0.246594
R953 VDD.n352 VDD.n351 0.246594
R954 VDD.n355 VDD.n354 0.246594
R955 VDD.n368 VDD.n367 0.246594
R956 VDD.n371 VDD.n370 0.246594
R957 VDD.n384 VDD.n383 0.246594
R958 VDD.n483 VDD.n482 0.239471
R959 VDD.n469 VDD.n468 0.239471
R960 VDD.n455 VDD.n454 0.239471
R961 VDD.n441 VDD.n440 0.239471
R962 VDD.n427 VDD.n426 0.239471
R963 VDD.n413 VDD.n412 0.239471
R964 VDD.n399 VDD.n398 0.239471
R965 VDD.n20 VDD.n19 0.232118
R966 VDD.n470 VDD.n28 0.232118
R967 VDD.n456 VDD.n36 0.232118
R968 VDD.n442 VDD.n44 0.232118
R969 VDD.n428 VDD.n52 0.232118
R970 VDD.n414 VDD.n60 0.232118
R971 VDD.n400 VDD.n68 0.232118
R972 VDD.n386 VDD.n76 0.232118
R973 VDD.n243 VDD.n240 0.229667
R974 VDD.n255 VDD.n254 0.229667
R975 VDD.n258 VDD.n234 0.229667
R976 VDD.n271 VDD.n270 0.229667
R977 VDD.n274 VDD.n228 0.229667
R978 VDD.n287 VDD.n286 0.229667
R979 VDD.n290 VDD.n222 0.229667
R980 VDD.n303 VDD.n302 0.229667
R981 VDD.n306 VDD.n216 0.229667
R982 VDD.n319 VDD.n318 0.229667
R983 VDD.n322 VDD.n210 0.229667
R984 VDD.n335 VDD.n334 0.229667
R985 VDD.n338 VDD.n204 0.229667
R986 VDD.n351 VDD.n350 0.229667
R987 VDD.n354 VDD.n198 0.229667
R988 VDD.n367 VDD.n366 0.229667
R989 VDD.n370 VDD.n192 0.229667
R990 VDD.n383 VDD.n382 0.229667
R991 VDD.n18 VDD.n17 0.124275
R992 VDD.n27 VDD.n23 0.124275
R993 VDD.n35 VDD.n31 0.124275
R994 VDD.n43 VDD.n39 0.124275
R995 VDD.n51 VDD.n47 0.124275
R996 VDD.n59 VDD.n55 0.124275
R997 VDD.n67 VDD.n63 0.124275
R998 VDD.n75 VDD.n71 0.124275
R999 VDD.n16 VDD.n3 0.121824
R1000 VDD.n481 VDD.n480 0.121824
R1001 VDD.n467 VDD.n466 0.121824
R1002 VDD.n453 VDD.n452 0.121824
R1003 VDD.n439 VDD.n438 0.121824
R1004 VDD.n425 VDD.n424 0.121824
R1005 VDD.n411 VDD.n410 0.121824
R1006 VDD.n397 VDD.n396 0.121824
R1007 VDD VDD.n20 0.113245
R1008 VDD.n470 VDD 0.113245
R1009 VDD.n456 VDD 0.113245
R1010 VDD.n442 VDD 0.113245
R1011 VDD.n428 VDD 0.113245
R1012 VDD.n414 VDD 0.113245
R1013 VDD.n400 VDD 0.113245
R1014 VDD.n386 VDD 0.113245
R1015 VDD.n117 VDD.n116 0.0804051
R1016 VDD.n127 VDD.n126 0.0804051
R1017 VDD.n137 VDD.n136 0.0804051
R1018 VDD.n147 VDD.n146 0.0804051
R1019 VDD.n157 VDD.n156 0.0804051
R1020 VDD.n167 VDD.n166 0.0804051
R1021 VDD.n177 VDD.n176 0.0804051
R1022 VDD.n187 VDD.n186 0.0804051
R1023 VDD VDD.n256 0.0708125
R1024 VDD VDD.n272 0.0708125
R1025 VDD VDD.n288 0.0708125
R1026 VDD VDD.n304 0.0708125
R1027 VDD VDD.n320 0.0708125
R1028 VDD VDD.n336 0.0708125
R1029 VDD VDD.n352 0.0708125
R1030 VDD VDD.n368 0.0708125
R1031 VDD VDD.n384 0.0708125
R1032 VDD.n17 VDD.n16 0.00295098
R1033 VDD.n480 VDD.n23 0.00295098
R1034 VDD.n466 VDD.n31 0.00295098
R1035 VDD.n452 VDD.n39 0.00295098
R1036 VDD.n438 VDD.n47 0.00295098
R1037 VDD.n424 VDD.n55 0.00295098
R1038 VDD.n410 VDD.n63 0.00295098
R1039 VDD.n396 VDD.n71 0.00295098
R1040 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 890.727
R1041 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 742.783
R1042 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 665.16
R1043 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 623.388
R1044 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 523.774
R1045 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 431.807
R1046 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 427.875
R1047 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 364.733
R1048 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 208.5
R1049 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 168.007
R1050 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R1051 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 31.2728
R1052 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R1053 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R1054 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R1055 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R1056 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 8.00471
R1057 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R1058 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R1059 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R1060 a_3116_2192.n3 a_3116_2192.n2 34.9195
R1061 a_3116_2192.n2 a_3116_2192.n0 25.5407
R1062 a_3116_2192.n2 a_3116_2192.n1 25.2907
R1063 a_3116_2192.n0 a_3116_2192.t5 5.8005
R1064 a_3116_2192.n0 a_3116_2192.t4 5.8005
R1065 a_3116_2192.n1 a_3116_2192.t3 5.8005
R1066 a_3116_2192.n1 a_3116_2192.t1 5.8005
R1067 a_3116_2192.n3 a_3116_2192.t2 5.8005
R1068 a_3116_2192.t0 a_3116_2192.n3 5.8005
R1069 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 879.481
R1070 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 742.783
R1071 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 665.16
R1072 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 623.388
R1073 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 523.774
R1074 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 431.807
R1075 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 427.875
R1076 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 357.26
R1077 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 208.537
R1078 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 168.077
R1079 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 75.5326
R1080 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R1081 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n7 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R1082 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 11.1806
R1083 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n7 10.5958
R1084 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R1085 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R1086 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 0.803118
R1087 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n7 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 0.23963
R1088 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 0.23963
R1089 VSS.n643 VSS.n77 6070.1
R1090 VSS.n458 VSS.n450 5774.44
R1091 VSS.n496 VSS.n311 5774.44
R1092 VSS.n346 VSS.n326 5774.44
R1093 VSS.n519 VSS.n228 5774.44
R1094 VSS.n263 VSS.n243 5774.44
R1095 VSS.n542 VSS.n194 5774.44
R1096 VSS.n473 VSS.n472 5774.44
R1097 VSS.n272 VSS.n200 4902.54
R1098 VSS.n278 VSS.n277 4902.54
R1099 VSS.n355 VSS.n283 4902.54
R1100 VSS.n361 VSS.n360 4902.54
R1101 VSS.n425 VSS.n366 4902.54
R1102 VSS.n441 VSS.n440 4902.54
R1103 VSS.n435 VSS.n434 4902.54
R1104 VSS.n550 VSS.n142 4200.9
R1105 VSS.n76 VSS.n75 4042.48
R1106 VSS.n397 VSS.n396 4042.48
R1107 VSS.n408 VSS.n407 4042.48
R1108 VSS.n310 VSS.n309 4042.48
R1109 VSS.n329 VSS.n328 4042.48
R1110 VSS.n227 VSS.n226 4042.48
R1111 VSS.n246 VSS.n245 4042.48
R1112 VSS.n156 VSS.n154 4042.48
R1113 VSS.n541 VSS.n200 3781.58
R1114 VSS.n277 VSS.n271 3781.58
R1115 VSS.n518 VSS.n283 3781.58
R1116 VSS.n360 VSS.n354 3781.58
R1117 VSS.n495 VSS.n366 3781.58
R1118 VSS.n449 VSS.n441 3781.58
R1119 VSS.n435 VSS.n405 3781.58
R1120 VSS.n399 VSS.n76 3140.17
R1121 VSS.n443 VSS.n397 3140.17
R1122 VSS.n415 VSS.n407 3140.17
R1123 VSS.n348 VSS.n310 3140.17
R1124 VSS.n336 VSS.n328 3140.17
R1125 VSS.n265 VSS.n227 3140.17
R1126 VSS.n253 VSS.n245 3140.17
R1127 VSS.n163 VSS.n156 3140.17
R1128 VSS.n652 VSS.n68 3120.05
R1129 VSS.n482 VSS.n389 3120.05
R1130 VSS.n378 VSS.n368 3120.05
R1131 VSS.n505 VSS.n302 3120.05
R1132 VSS.n295 VSS.n285 3120.05
R1133 VSS.n528 VSS.n219 3120.05
R1134 VSS.n212 VSS.n202 3120.05
R1135 VSS.n544 VSS.n144 3120.05
R1136 VSS.n195 VSS.n141 2421.55
R1137 VSS.n652 VSS.n67 2350.81
R1138 VSS.n482 VSS.n388 2350.81
R1139 VSS.n493 VSS.n368 2350.81
R1140 VSS.n505 VSS.n301 2350.81
R1141 VSS.n516 VSS.n285 2350.81
R1142 VSS.n528 VSS.n218 2350.81
R1143 VSS.n539 VSS.n202 2350.81
R1144 VSS.n548 VSS.n144 2350.81
R1145 VSS.n184 VSS.n180 2235.89
R1146 VSS.n236 VSS.n3 2235.89
R1147 VSS.n234 VSS.n12 2235.89
R1148 VSS.n319 VSS.n21 2235.89
R1149 VSS.n317 VSS.n30 2235.89
R1150 VSS.n451 VSS.n39 2235.89
R1151 VSS.n459 VSS.n48 2235.89
R1152 VSS.n470 VSS.n57 2235.89
R1153 VSS.n192 VSS.n172 2230.09
R1154 VSS.n239 VSS.n5 2230.09
R1155 VSS.n230 VSS.n14 2230.09
R1156 VSS.n322 VSS.n23 2230.09
R1157 VSS.n313 VSS.n32 2230.09
R1158 VSS.n454 VSS.n41 2230.09
R1159 VSS.n462 VSS.n50 2230.09
R1160 VSS.n466 VSS.n59 2230.09
R1161 VSS.n641 VSS.n78 2120.77
R1162 VSS.n433 VSS.n78 2120.77
R1163 VSS.n437 VSS.n436 2120.77
R1164 VSS.n436 VSS.n91 2120.77
R1165 VSS.n428 VSS.n427 2120.77
R1166 VSS.n427 VSS.n98 2120.77
R1167 VSS.n364 VSS.n363 2120.77
R1168 VSS.n363 VSS.n105 2120.77
R1169 VSS.n358 VSS.n357 2120.77
R1170 VSS.n357 VSS.n112 2120.77
R1171 VSS.n281 VSS.n280 2120.77
R1172 VSS.n280 VSS.n119 2120.77
R1173 VSS.n275 VSS.n274 2120.77
R1174 VSS.n274 VSS.n126 2120.77
R1175 VSS.n198 VSS.n197 2120.77
R1176 VSS.n197 VSS.n133 2120.77
R1177 VSS.n140 VSS.n136 2120.77
R1178 VSS.n553 VSS.n140 2120.77
R1179 VSS.n646 VSS.n76 1915.82
R1180 VSS.n476 VSS.n397 1915.82
R1181 VSS.n422 VSS.n407 1915.82
R1182 VSS.n499 VSS.n310 1915.82
R1183 VSS.n343 VSS.n328 1915.82
R1184 VSS.n522 VSS.n227 1915.82
R1185 VSS.n260 VSS.n245 1915.82
R1186 VSS.n170 VSS.n156 1915.82
R1187 VSS.n646 VSS.n71 1832.1
R1188 VSS.n476 VSS.n392 1832.1
R1189 VSS.n422 VSS.n409 1832.1
R1190 VSS.n499 VSS.n305 1832.1
R1191 VSS.n343 VSS.n330 1832.1
R1192 VSS.n522 VSS.n222 1832.1
R1193 VSS.n260 VSS.n247 1832.1
R1194 VSS.n170 VSS.n157 1832.1
R1195 VSS.n200 VSS.n199 1630.46
R1196 VSS.n277 VSS.n276 1630.46
R1197 VSS.n283 VSS.n282 1630.46
R1198 VSS.n360 VSS.n359 1630.46
R1199 VSS.n366 VSS.n365 1630.46
R1200 VSS.n441 VSS.n429 1630.46
R1201 VSS.n438 VSS.n435 1630.46
R1202 VSS.n402 VSS.n67 1562.99
R1203 VSS.n446 VSS.n388 1562.99
R1204 VSS.n493 VSS.n367 1562.99
R1205 VSS.n351 VSS.n301 1562.99
R1206 VSS.n516 VSS.n284 1562.99
R1207 VSS.n268 VSS.n218 1562.99
R1208 VSS.n539 VSS.n201 1562.99
R1209 VSS.n548 VSS.n143 1562.99
R1210 VSS.n181 VSS.n172 1411.83
R1211 VSS.n240 VSS.n239 1411.83
R1212 VSS.n231 VSS.n230 1411.83
R1213 VSS.n323 VSS.n322 1411.83
R1214 VSS.n314 VSS.n313 1411.83
R1215 VSS.n455 VSS.n454 1411.83
R1216 VSS.n463 VSS.n462 1411.83
R1217 VSS.n467 VSS.n466 1411.83
R1218 VSS.n550 VSS.n549 1255.49
R1219 VSS.n650 VSS.n70 1226.74
R1220 VSS.n480 VSS.n391 1226.74
R1221 VSS.n418 VSS.n412 1226.74
R1222 VSS.n503 VSS.n304 1226.74
R1223 VSS.n339 VSS.n333 1226.74
R1224 VSS.n526 VSS.n221 1226.74
R1225 VSS.n256 VSS.n250 1226.74
R1226 VSS.n166 VSS.n160 1226.74
R1227 VSS.n75 VSS.n71 1068.72
R1228 VSS.n396 VSS.n392 1068.72
R1229 VSS.n409 VSS.n408 1068.72
R1230 VSS.n309 VSS.n305 1068.72
R1231 VSS.n330 VSS.n329 1068.72
R1232 VSS.n226 VSS.n222 1068.72
R1233 VSS.n247 VSS.n246 1068.72
R1234 VSS.n157 VSS.n154 1068.72
R1235 VSS.t257 VSS.n460 994.611
R1236 VSS.t61 VSS.n452 994.611
R1237 VSS.n318 VSS.t209 994.611
R1238 VSS.t63 VSS.n320 994.611
R1239 VSS.n235 VSS.t338 994.611
R1240 VSS.t324 VSS.n237 994.611
R1241 VSS.t262 VSS.n142 994.611
R1242 VSS.n471 VSS.t30 994.611
R1243 VSS.t276 VSS.n464 955.091
R1244 VSS.n465 VSS.t226 955.091
R1245 VSS.t73 VSS.n456 955.091
R1246 VSS.n457 VSS.t249 955.091
R1247 VSS.n315 VSS.t332 955.091
R1248 VSS.t284 VSS.n312 955.091
R1249 VSS.t150 VSS.n324 955.091
R1250 VSS.n325 VSS.t176 955.091
R1251 VSS.n232 VSS.t194 955.091
R1252 VSS.t201 VSS.n229 955.091
R1253 VSS.t278 VSS.n241 955.091
R1254 VSS.n242 VSS.t296 955.091
R1255 VSS.n182 VSS.t334 955.091
R1256 VSS.n193 VSS.t303 955.091
R1257 VSS.n468 VSS.t370 955.091
R1258 VSS.t343 VSS.n77 955.091
R1259 VSS.n461 VSS.t353 935.33
R1260 VSS.n453 VSS.t131 935.33
R1261 VSS.t100 VSS.n316 935.33
R1262 VSS.n321 VSS.t204 935.33
R1263 VSS.t322 VSS.n233 935.33
R1264 VSS.n238 VSS.t169 935.33
R1265 VSS.n183 VSS.t22 935.33
R1266 VSS.t197 VSS.n469 935.33
R1267 VSS.n644 VSS.n643 886.567
R1268 VSS.n543 VSS.n542 832.486
R1269 VSS.n263 VSS.n262 832.486
R1270 VSS.n520 VSS.n519 832.486
R1271 VSS.n346 VSS.n345 832.486
R1272 VSS.n497 VSS.n496 832.486
R1273 VSS.n450 VSS.n424 832.486
R1274 VSS.n474 VSS.n473 832.486
R1275 VSS.t388 VSS.n195 815.229
R1276 VSS.n196 VSS.t24 815.229
R1277 VSS.t159 VSS.n196 815.229
R1278 VSS.n199 VSS.t80 815.229
R1279 VSS.t8 VSS.n272 815.229
R1280 VSS.n273 VSS.t146 815.229
R1281 VSS.t156 VSS.n273 815.229
R1282 VSS.n276 VSS.t47 815.229
R1283 VSS.t267 VSS.n278 815.229
R1284 VSS.n279 VSS.t372 815.229
R1285 VSS.t231 VSS.n279 815.229
R1286 VSS.n282 VSS.t239 815.229
R1287 VSS.t143 VSS.n355 815.229
R1288 VSS.n356 VSS.t286 815.229
R1289 VSS.t328 VSS.n356 815.229
R1290 VSS.n359 VSS.t365 815.229
R1291 VSS.t247 VSS.n361 815.229
R1292 VSS.n362 VSS.t349 815.229
R1293 VSS.t115 VSS.n362 815.229
R1294 VSS.n365 VSS.t394 815.229
R1295 VSS.t123 VSS.n425 815.229
R1296 VSS.n426 VSS.t121 815.229
R1297 VSS.t2 VSS.n426 815.229
R1298 VSS.n429 VSS.t0 815.229
R1299 VSS.n440 VSS.t107 815.229
R1300 VSS.t112 VSS.n439 815.229
R1301 VSS.n439 VSS.t318 815.229
R1302 VSS.t315 VSS.n438 815.229
R1303 VSS.n434 VSS.t313 815.229
R1304 VSS.t307 VSS.n432 815.229
R1305 VSS.n432 VSS.t171 815.229
R1306 VSS.n399 VSS.n70 742.855
R1307 VSS.n443 VSS.n391 742.855
R1308 VSS.n415 VSS.n412 742.855
R1309 VSS.n348 VSS.n304 742.855
R1310 VSS.n336 VSS.n333 742.855
R1311 VSS.n265 VSS.n221 742.855
R1312 VSS.n253 VSS.n250 742.855
R1313 VSS.n163 VSS.n160 742.855
R1314 VSS.n472 VSS.n465 605.989
R1315 VSS.n458 VSS.n457 605.989
R1316 VSS.n312 VSS.n311 605.989
R1317 VSS.n326 VSS.n325 605.989
R1318 VSS.n229 VSS.n228 605.989
R1319 VSS.n243 VSS.n242 605.989
R1320 VSS.n194 VSS.n193 605.989
R1321 VSS.n460 VSS.n458 592.814
R1322 VSS.n452 VSS.n311 592.814
R1323 VSS.n326 VSS.n318 592.814
R1324 VSS.n320 VSS.n228 592.814
R1325 VSS.n243 VSS.n235 592.814
R1326 VSS.n237 VSS.n194 592.814
R1327 VSS.n472 VSS.n471 592.814
R1328 VSS.t90 VSS.t257 579.641
R1329 VSS.t224 VSS.t90 579.641
R1330 VSS.t353 VSS.t224 579.641
R1331 VSS.t259 VSS.t276 579.641
R1332 VSS.t78 VSS.t259 579.641
R1333 VSS.t226 VSS.t78 579.641
R1334 VSS.t190 VSS.t61 579.641
R1335 VSS.t381 VSS.t190 579.641
R1336 VSS.t131 VSS.t381 579.641
R1337 VSS.t158 VSS.t73 579.641
R1338 VSS.t288 VSS.t158 579.641
R1339 VSS.t249 VSS.t288 579.641
R1340 VSS.t209 VSS.t211 579.641
R1341 VSS.t211 VSS.t236 579.641
R1342 VSS.t236 VSS.t100 579.641
R1343 VSS.t332 VSS.t206 579.641
R1344 VSS.t206 VSS.t188 579.641
R1345 VSS.t188 VSS.t284 579.641
R1346 VSS.t152 VSS.t63 579.641
R1347 VSS.t355 VSS.t152 579.641
R1348 VSS.t204 VSS.t355 579.641
R1349 VSS.t173 VSS.t150 579.641
R1350 VSS.t16 VSS.t173 579.641
R1351 VSS.t176 VSS.t16 579.641
R1352 VSS.t338 VSS.t280 579.641
R1353 VSS.t280 VSS.t75 579.641
R1354 VSS.t75 VSS.t322 579.641
R1355 VSS.t194 VSS.t356 579.641
R1356 VSS.t356 VSS.t186 579.641
R1357 VSS.t186 VSS.t201 579.641
R1358 VSS.t14 VSS.t324 579.641
R1359 VSS.t299 VSS.t14 579.641
R1360 VSS.t169 VSS.t299 579.641
R1361 VSS.t66 VSS.t278 579.641
R1362 VSS.t234 VSS.t66 579.641
R1363 VSS.t296 VSS.t234 579.641
R1364 VSS.t260 VSS.t262 579.641
R1365 VSS.t306 VSS.t260 579.641
R1366 VSS.t22 VSS.t306 579.641
R1367 VSS.t334 VSS.t264 579.641
R1368 VSS.t264 VSS.t330 579.641
R1369 VSS.t330 VSS.t303 579.641
R1370 VSS.t30 VSS.t68 579.641
R1371 VSS.t68 VSS.t340 579.641
R1372 VSS.t340 VSS.t197 579.641
R1373 VSS.t370 VSS.t67 579.641
R1374 VSS.t67 VSS.t70 579.641
R1375 VSS.t70 VSS.t343 579.641
R1376 VSS.t222 VSS.t388 491.372
R1377 VSS.t351 VSS.t222 491.372
R1378 VSS.t24 VSS.t351 491.372
R1379 VSS.t213 VSS.t377 491.372
R1380 VSS.t80 VSS.t213 491.372
R1381 VSS.t336 VSS.t8 491.372
R1382 VSS.t94 VSS.t336 491.372
R1383 VSS.t146 VSS.t94 491.372
R1384 VSS.t346 VSS.t26 491.372
R1385 VSS.t47 VSS.t346 491.372
R1386 VSS.t44 VSS.t267 491.372
R1387 VSS.t245 VSS.t44 491.372
R1388 VSS.t372 VSS.t245 491.372
R1389 VSS.t199 VSS.t229 491.372
R1390 VSS.t239 VSS.t199 491.372
R1391 VSS.t390 VSS.t143 491.372
R1392 VSS.t207 VSS.t390 491.372
R1393 VSS.t286 VSS.t207 491.372
R1394 VSS.t368 VSS.t97 491.372
R1395 VSS.t365 VSS.t368 491.372
R1396 VSS.t163 VSS.t247 491.372
R1397 VSS.t237 VSS.t163 491.372
R1398 VSS.t349 VSS.t237 491.372
R1399 VSS.t398 VSS.t294 491.372
R1400 VSS.t394 VSS.t398 491.372
R1401 VSS.t119 VSS.t123 491.372
R1402 VSS.t125 VSS.t119 491.372
R1403 VSS.t121 VSS.t125 491.372
R1404 VSS.t18 VSS.t5 491.372
R1405 VSS.t0 VSS.t18 491.372
R1406 VSS.t107 VSS.t110 491.372
R1407 VSS.t110 VSS.t104 491.372
R1408 VSS.t104 VSS.t112 491.372
R1409 VSS.t320 VSS.t251 491.372
R1410 VSS.t251 VSS.t315 491.372
R1411 VSS.t313 VSS.t309 491.372
R1412 VSS.t309 VSS.t311 491.372
R1413 VSS.t311 VSS.t307 491.372
R1414 VSS.t377 VSS.t159 477.411
R1415 VSS.t26 VSS.t156 477.411
R1416 VSS.t229 VSS.t231 477.411
R1417 VSS.t97 VSS.t328 477.411
R1418 VSS.t294 VSS.t115 477.411
R1419 VSS.t5 VSS.t2 477.411
R1420 VSS.t318 VSS.t320 477.411
R1421 VSS.t171 VSS.t292 471.786
R1422 VSS.n553 VSS.t265 463.868
R1423 VSS.n541 VSS.n540 446.182
R1424 VSS.n271 VSS.n270 446.182
R1425 VSS.n518 VSS.n517 446.182
R1426 VSS.n354 VSS.n353 446.182
R1427 VSS.n495 VSS.n494 446.182
R1428 VSS.n449 VSS.n448 446.182
R1429 VSS.n405 VSS.n404 446.182
R1430 VSS.n643 VSS.n642 441.358
R1431 VSS.n542 VSS.n541 413.346
R1432 VSS.n271 VSS.n263 413.346
R1433 VSS.n519 VSS.n518 413.346
R1434 VSS.n354 VSS.n346 413.346
R1435 VSS.n496 VSS.n495 413.346
R1436 VSS.n450 VSS.n449 413.346
R1437 VSS.n473 VSS.n405 413.346
R1438 VSS.n402 VSS.n70 356.277
R1439 VSS.n446 VSS.n391 356.277
R1440 VSS.n412 VSS.n367 356.277
R1441 VSS.n351 VSS.n304 356.277
R1442 VSS.n333 VSS.n284 356.277
R1443 VSS.n268 VSS.n221 356.277
R1444 VSS.n250 VSS.n201 356.277
R1445 VSS.n160 VSS.n143 356.277
R1446 VSS.t76 VSS.n552 346.868
R1447 VSS.n552 VSS.t379 346.868
R1448 VSS.n642 VSS.t290 346.868
R1449 VSS.n549 VSS.t384 338.017
R1450 VSS.n543 VSS.t103 338.017
R1451 VSS.n540 VSS.t32 338.017
R1452 VSS.n262 VSS.t166 338.017
R1453 VSS.n270 VSS.t59 338.017
R1454 VSS.t65 VSS.n520 338.017
R1455 VSS.n517 VSS.t51 338.017
R1456 VSS.n345 VSS.t145 338.017
R1457 VSS.n353 VSS.t326 338.017
R1458 VSS.t298 VSS.n497 338.017
R1459 VSS.n494 VSS.t129 338.017
R1460 VSS.n424 VSS.t165 338.017
R1461 VSS.n448 VSS.t141 338.017
R1462 VSS.t221 VSS.n474 338.017
R1463 VSS.n404 VSS.t382 338.017
R1464 VSS.t114 VSS.n644 338.017
R1465 VSS.n550 VSS.n141 301.728
R1466 VSS.n75 VSS.n68 281.135
R1467 VSS.n396 VSS.n389 281.135
R1468 VSS.n408 VSS.n378 281.135
R1469 VSS.n309 VSS.n302 281.135
R1470 VSS.n329 VSS.n295 281.135
R1471 VSS.n226 VSS.n219 281.135
R1472 VSS.n246 VSS.n212 281.135
R1473 VSS.n544 VSS.n154 281.135
R1474 VSS.n248 VSS.n211 262.659
R1475 VSS.n225 VSS.n224 262.659
R1476 VSS.n331 VSS.n294 262.659
R1477 VSS.n308 VSS.n307 262.659
R1478 VSS.n410 VSS.n377 262.659
R1479 VSS.n395 VSS.n394 262.659
R1480 VSS.n74 VSS.n73 262.659
R1481 VSS.n158 VSS.n152 262.659
R1482 VSS.t265 VSS.t154 209.071
R1483 VSS.t154 VSS.t282 209.071
R1484 VSS.t282 VSS.t76 209.071
R1485 VSS.t379 VSS.t28 209.071
R1486 VSS.t28 VSS.t272 209.071
R1487 VSS.t272 VSS.t40 209.071
R1488 VSS.t292 VSS.t301 209.071
R1489 VSS.t301 VSS.t290 209.071
R1490 VSS.n252 VSS.n248 204.031
R1491 VSS.n264 VSS.n225 204.031
R1492 VSS.n335 VSS.n331 204.031
R1493 VSS.n347 VSS.n308 204.031
R1494 VSS.n414 VSS.n410 204.031
R1495 VSS.n442 VSS.n395 204.031
R1496 VSS.n398 VSS.n74 204.031
R1497 VSS.n162 VSS.n158 204.031
R1498 VSS.n537 VSS.n536 202.725
R1499 VSS.n529 VSS.n217 202.725
R1500 VSS.n514 VSS.n513 202.725
R1501 VSS.n506 VSS.n300 202.725
R1502 VSS.n491 VSS.n490 202.725
R1503 VSS.n483 VSS.n387 202.725
R1504 VSS.n653 VSS.n63 202.725
R1505 VSS.n546 VSS.n545 202.725
R1506 VSS.t361 VSS.t53 169.975
R1507 VSS.t392 VSS.t357 169.975
R1508 VSS.t180 VSS.t392 169.975
R1509 VSS.t93 VSS.t180 169.975
R1510 VSS.t228 VSS.t93 169.975
R1511 VSS.t184 VSS.t228 169.975
R1512 VSS.t168 VSS.t193 169.975
R1513 VSS.t305 VSS.t168 169.975
R1514 VSS.t103 VSS.t305 169.975
R1515 VSS.t55 VSS.t255 169.975
R1516 VSS.t359 VSS.t363 169.975
R1517 VSS.t11 VSS.t359 169.975
R1518 VSS.t128 VSS.t11 169.975
R1519 VSS.t203 VSS.t128 169.975
R1520 VSS.t376 VSS.t203 169.975
R1521 VSS.t178 VSS.t134 169.975
R1522 VSS.t118 VSS.t178 169.975
R1523 VSS.t166 VSS.t118 169.975
R1524 VSS.t34 VSS.t139 169.975
R1525 VSS.t88 VSS.t386 169.975
R1526 VSS.t386 VSS.t271 169.975
R1527 VSS.t10 VSS.t271 169.975
R1528 VSS.t10 VSS.t196 169.975
R1529 VSS.t196 VSS.t174 169.975
R1530 VSS.t92 VSS.t161 169.975
R1531 VSS.t161 VSS.t127 169.975
R1532 VSS.t127 VSS.t65 169.975
R1533 VSS.t135 VSS.t215 169.975
R1534 VSS.t49 VSS.t243 169.975
R1535 VSS.t300 VSS.t49 169.975
R1536 VSS.t179 VSS.t300 169.975
R1537 VSS.t374 VSS.t179 169.975
R1538 VSS.t46 VSS.t374 169.975
R1539 VSS.t269 VSS.t133 169.975
R1540 VSS.t270 VSS.t269 169.975
R1541 VSS.t145 VSS.t270 169.975
R1542 VSS.t217 VSS.t137 169.975
R1543 VSS.t341 VSS.t57 169.975
R1544 VSS.t57 VSS.t99 169.975
R1545 VSS.t175 VSS.t99 169.975
R1546 VSS.t175 VSS.t102 169.975
R1547 VSS.t102 VSS.t233 169.975
R1548 VSS.t43 VSS.t367 169.975
R1549 VSS.t367 VSS.t72 169.975
R1550 VSS.t72 VSS.t298 169.975
R1551 VSS.t86 VSS.t241 169.975
R1552 VSS.t219 VSS.t82 169.975
R1553 VSS.t348 VSS.t219 169.975
R1554 VSS.t162 VSS.t348 169.975
R1555 VSS.t185 VSS.t162 169.975
R1556 VSS.t167 VSS.t185 169.975
R1557 VSS.t397 VSS.t396 169.975
R1558 VSS.t181 VSS.t397 169.975
R1559 VSS.t165 VSS.t181 169.975
R1560 VSS.t148 VSS.t36 169.975
R1561 VSS.t253 VSS.t84 169.975
R1562 VSS.t84 VSS.t21 169.975
R1563 VSS.t7 VSS.t21 169.975
R1564 VSS.t7 VSS.t117 169.975
R1565 VSS.t117 VSS.t345 169.975
R1566 VSS.t20 VSS.t4 169.975
R1567 VSS.t4 VSS.t225 169.975
R1568 VSS.t225 VSS.t221 169.975
R1569 VSS.t12 VSS.t182 169.975
R1570 VSS.t38 VSS.t274 169.975
R1571 VSS.t274 VSS.t96 169.975
R1572 VSS.t42 VSS.t96 169.975
R1573 VSS.t42 VSS.t106 169.975
R1574 VSS.t106 VSS.t192 169.975
R1575 VSS.t317 VSS.t375 169.975
R1576 VSS.t375 VSS.t109 169.975
R1577 VSS.t109 VSS.t114 169.975
R1578 VSS.n164 VSS.t361 168.042
R1579 VSS.n254 VSS.t55 168.042
R1580 VSS.t139 VSS.n266 168.042
R1581 VSS.n337 VSS.t135 168.042
R1582 VSS.t137 VSS.n349 168.042
R1583 VSS.n416 VSS.t86 168.042
R1584 VSS.t36 VSS.n444 168.042
R1585 VSS.t182 VSS.n400 168.042
R1586 VSS.n538 VSS.n537 152.744
R1587 VSS.n529 VSS.n213 152.744
R1588 VSS.n515 VSS.n514 152.744
R1589 VSS.n506 VSS.n296 152.744
R1590 VSS.n492 VSS.n491 152.744
R1591 VSS.n483 VSS.n379 152.744
R1592 VSS.n653 VSS.n66 152.744
R1593 VSS.n547 VSS.n546 152.744
R1594 VSS.n185 VSS.n179 138.52
R1595 VSS.n708 VSS.n0 138.52
R1596 VSS.n700 VSS.n9 138.52
R1597 VSS.n692 VSS.n18 138.52
R1598 VSS.n684 VSS.n27 138.52
R1599 VSS.n676 VSS.n36 138.52
R1600 VSS.n668 VSS.n45 138.52
R1601 VSS.n660 VSS.n54 138.52
R1602 VSS.n191 VSS.n173 138.144
R1603 VSS.n707 VSS.n706 138.144
R1604 VSS.n699 VSS.n698 138.144
R1605 VSS.n691 VSS.n690 138.144
R1606 VSS.n683 VSS.n682 138.144
R1607 VSS.n675 VSS.n674 138.144
R1608 VSS.n667 VSS.n666 138.144
R1609 VSS.n659 VSS.n658 138.144
R1610 VSS.n567 VSS.n566 137.46
R1611 VSS.n577 VSS.n576 137.46
R1612 VSS.n587 VSS.n586 137.46
R1613 VSS.n597 VSS.n596 137.46
R1614 VSS.n607 VSS.n606 137.46
R1615 VSS.n617 VSS.n616 137.46
R1616 VSS.n627 VSS.n626 137.46
R1617 VSS.n430 VSS.n84 137.46
R1618 VSS.n554 VSS.n137 137.46
R1619 VSS.n568 VSS.n127 136.661
R1620 VSS.n578 VSS.n120 136.661
R1621 VSS.n588 VSS.n113 136.661
R1622 VSS.n598 VSS.n106 136.661
R1623 VSS.n608 VSS.n99 136.661
R1624 VSS.n618 VSS.n92 136.661
R1625 VSS.n628 VSS.n85 136.661
R1626 VSS.n640 VSS.n79 136.661
R1627 VSS.n561 VSS.n560 136.661
R1628 VSS.n259 VSS.n248 124.481
R1629 VSS.n523 VSS.n225 124.481
R1630 VSS.n342 VSS.n331 124.481
R1631 VSS.n500 VSS.n308 124.481
R1632 VSS.n421 VSS.n410 124.481
R1633 VSS.n477 VSS.n395 124.481
R1634 VSS.n647 VSS.n74 124.481
R1635 VSS.n169 VSS.n158 124.481
R1636 VSS.n259 VSS.n258 119.04
R1637 VSS.n524 VSS.n523 119.04
R1638 VSS.n342 VSS.n341 119.04
R1639 VSS.n501 VSS.n500 119.04
R1640 VSS.n421 VSS.n420 119.04
R1641 VSS.n478 VSS.n477 119.04
R1642 VSS.n648 VSS.n647 119.04
R1643 VSS.n169 VSS.n168 119.04
R1644 VSS.n566 VSS.n133 117.338
R1645 VSS.n198 VSS.n127 117.338
R1646 VSS.n576 VSS.n126 117.338
R1647 VSS.n275 VSS.n120 117.338
R1648 VSS.n586 VSS.n119 117.338
R1649 VSS.n281 VSS.n113 117.338
R1650 VSS.n596 VSS.n112 117.338
R1651 VSS.n358 VSS.n106 117.338
R1652 VSS.n606 VSS.n105 117.338
R1653 VSS.n364 VSS.n99 117.338
R1654 VSS.n616 VSS.n98 117.338
R1655 VSS.n428 VSS.n92 117.338
R1656 VSS.n626 VSS.n91 117.338
R1657 VSS.n437 VSS.n85 117.338
R1658 VSS.n433 VSS.n84 117.338
R1659 VSS.n641 VSS.n640 117.338
R1660 VSS.n561 VSS.n136 117.338
R1661 VSS.n554 VSS.n553 117.338
R1662 VSS.n141 VSS.n136 117.001
R1663 VSS.n195 VSS.n133 117.001
R1664 VSS.n199 VSS.n198 117.001
R1665 VSS.n272 VSS.n126 117.001
R1666 VSS.n276 VSS.n275 117.001
R1667 VSS.n278 VSS.n119 117.001
R1668 VSS.n282 VSS.n281 117.001
R1669 VSS.n355 VSS.n112 117.001
R1670 VSS.n359 VSS.n358 117.001
R1671 VSS.n361 VSS.n105 117.001
R1672 VSS.n365 VSS.n364 117.001
R1673 VSS.n425 VSS.n98 117.001
R1674 VSS.n429 VSS.n428 117.001
R1675 VSS.n440 VSS.n91 117.001
R1676 VSS.n438 VSS.n437 117.001
R1677 VSS.n434 VSS.n433 117.001
R1678 VSS.n642 VSS.n641 117.001
R1679 VSS.n145 VSS.n143 117.001
R1680 VSS.n161 VSS.n143 117.001
R1681 VSS.n203 VSS.n201 117.001
R1682 VSS.n251 VSS.n201 117.001
R1683 VSS.n268 VSS.n267 117.001
R1684 VSS.n269 VSS.n268 117.001
R1685 VSS.n286 VSS.n284 117.001
R1686 VSS.n334 VSS.n284 117.001
R1687 VSS.n351 VSS.n350 117.001
R1688 VSS.n352 VSS.n351 117.001
R1689 VSS.n369 VSS.n367 117.001
R1690 VSS.n413 VSS.n367 117.001
R1691 VSS.n446 VSS.n445 117.001
R1692 VSS.n447 VSS.n446 117.001
R1693 VSS.n402 VSS.n401 117.001
R1694 VSS.n403 VSS.n402 117.001
R1695 VSS.n192 VSS.n191 104.257
R1696 VSS.n180 VSS.n179 104.257
R1697 VSS.n706 VSS.n5 104.257
R1698 VSS.n236 VSS.n0 104.257
R1699 VSS.n698 VSS.n14 104.257
R1700 VSS.n234 VSS.n9 104.257
R1701 VSS.n690 VSS.n23 104.257
R1702 VSS.n319 VSS.n18 104.257
R1703 VSS.n682 VSS.n32 104.257
R1704 VSS.n317 VSS.n27 104.257
R1705 VSS.n674 VSS.n41 104.257
R1706 VSS.n451 VSS.n36 104.257
R1707 VSS.n666 VSS.n50 104.257
R1708 VSS.n459 VSS.n45 104.257
R1709 VSS.n470 VSS.n54 104.257
R1710 VSS.n658 VSS.n59 104.257
R1711 VSS.n538 VSS.n203 101.555
R1712 VSS.n267 VSS.n213 101.555
R1713 VSS.n515 VSS.n286 101.555
R1714 VSS.n350 VSS.n296 101.555
R1715 VSS.n492 VSS.n369 101.555
R1716 VSS.n445 VSS.n379 101.555
R1717 VSS.n401 VSS.n66 101.555
R1718 VSS.n547 VSS.n145 101.555
R1719 VSS.n460 VSS.n459 97.5005
R1720 VSS.n465 VSS.n50 97.5005
R1721 VSS.n452 VSS.n451 97.5005
R1722 VSS.n457 VSS.n41 97.5005
R1723 VSS.n318 VSS.n317 97.5005
R1724 VSS.n312 VSS.n32 97.5005
R1725 VSS.n320 VSS.n319 97.5005
R1726 VSS.n325 VSS.n23 97.5005
R1727 VSS.n235 VSS.n234 97.5005
R1728 VSS.n229 VSS.n14 97.5005
R1729 VSS.n237 VSS.n236 97.5005
R1730 VSS.n242 VSS.n5 97.5005
R1731 VSS.n180 VSS.n142 97.5005
R1732 VSS.n193 VSS.n192 97.5005
R1733 VSS.n471 VSS.n470 97.5005
R1734 VSS.n77 VSS.n59 97.5005
R1735 VSS.n181 VSS.n175 92.3255
R1736 VSS.n240 VSS.n4 92.3255
R1737 VSS.n231 VSS.n13 92.3255
R1738 VSS.n323 VSS.n22 92.3255
R1739 VSS.n314 VSS.n31 92.3255
R1740 VSS.n455 VSS.n40 92.3255
R1741 VSS.n463 VSS.n49 92.3255
R1742 VSS.n467 VSS.n58 92.3255
R1743 VSS.n161 VSS.t384 86.9189
R1744 VSS.n251 VSS.t32 86.9189
R1745 VSS.t59 VSS.n269 86.9189
R1746 VSS.n334 VSS.t51 86.9189
R1747 VSS.t326 VSS.n352 86.9189
R1748 VSS.n413 VSS.t129 86.9189
R1749 VSS.t141 VSS.n447 86.9189
R1750 VSS.t382 VSS.n403 86.9189
R1751 VSS.n176 VSS.t23 84.5161
R1752 VSS.n188 VSS.t335 84.5161
R1753 VSS.n710 VSS.t170 84.5161
R1754 VSS.n7 VSS.t279 84.5161
R1755 VSS.n702 VSS.t323 84.5161
R1756 VSS.n16 VSS.t195 84.5161
R1757 VSS.n694 VSS.t205 84.5161
R1758 VSS.n25 VSS.t151 84.5161
R1759 VSS.n686 VSS.t101 84.5161
R1760 VSS.n34 VSS.t333 84.5161
R1761 VSS.n678 VSS.t132 84.5161
R1762 VSS.n43 VSS.t74 84.5161
R1763 VSS.n670 VSS.t354 84.5161
R1764 VSS.n52 VSS.t277 84.5161
R1765 VSS.n662 VSS.t198 84.5161
R1766 VSS.n61 VSS.t371 84.5161
R1767 VSS.t53 VSS.n161 83.0558
R1768 VSS.t193 VSS.n171 83.0558
R1769 VSS.t255 VSS.n251 83.0558
R1770 VSS.t134 VSS.n261 83.0558
R1771 VSS.n269 VSS.t34 83.0558
R1772 VSS.n521 VSS.t92 83.0558
R1773 VSS.t215 VSS.n334 83.0558
R1774 VSS.t133 VSS.n344 83.0558
R1775 VSS.n352 VSS.t217 83.0558
R1776 VSS.n498 VSS.t43 83.0558
R1777 VSS.t241 VSS.n413 83.0558
R1778 VSS.t396 VSS.n423 83.0558
R1779 VSS.n447 VSS.t148 83.0558
R1780 VSS.n475 VSS.t20 83.0558
R1781 VSS.n403 VSS.t12 83.0558
R1782 VSS.n645 VSS.t317 83.0558
R1783 VSS.n257 VSS.n249 79.7072
R1784 VSS.n525 VSS.n223 79.7072
R1785 VSS.n340 VSS.n332 79.7072
R1786 VSS.n502 VSS.n306 79.7072
R1787 VSS.n419 VSS.n411 79.7072
R1788 VSS.n479 VSS.n393 79.7072
R1789 VSS.n649 VSS.n72 79.7072
R1790 VSS.n167 VSS.n159 79.7072
R1791 VSS.n464 VSS.n463 73.1255
R1792 VSS.n456 VSS.n455 73.1255
R1793 VSS.n315 VSS.n314 73.1255
R1794 VSS.n324 VSS.n323 73.1255
R1795 VSS.n232 VSS.n231 73.1255
R1796 VSS.n241 VSS.n240 73.1255
R1797 VSS.n182 VSS.n181 73.1255
R1798 VSS.n163 VSS.n162 73.1255
R1799 VSS.n164 VSS.n163 73.1255
R1800 VSS.n253 VSS.n252 73.1255
R1801 VSS.n254 VSS.n253 73.1255
R1802 VSS.n265 VSS.n264 73.1255
R1803 VSS.n266 VSS.n265 73.1255
R1804 VSS.n336 VSS.n335 73.1255
R1805 VSS.n337 VSS.n336 73.1255
R1806 VSS.n348 VSS.n347 73.1255
R1807 VSS.n349 VSS.n348 73.1255
R1808 VSS.n415 VSS.n414 73.1255
R1809 VSS.n416 VSS.n415 73.1255
R1810 VSS.n443 VSS.n442 73.1255
R1811 VSS.n444 VSS.n443 73.1255
R1812 VSS.n399 VSS.n398 73.1255
R1813 VSS.n400 VSS.n399 73.1255
R1814 VSS.n468 VSS.n467 73.1255
R1815 VSS.n175 VSS.n173 72.5338
R1816 VSS.n707 VSS.n4 72.5338
R1817 VSS.n699 VSS.n13 72.5338
R1818 VSS.n691 VSS.n22 72.5338
R1819 VSS.n683 VSS.n31 72.5338
R1820 VSS.n675 VSS.n40 72.5338
R1821 VSS.n667 VSS.n49 72.5338
R1822 VSS.n659 VSS.n58 72.5338
R1823 VSS.n258 VSS.n211 69.4405
R1824 VSS.n524 VSS.n224 69.4405
R1825 VSS.n341 VSS.n294 69.4405
R1826 VSS.n501 VSS.n307 69.4405
R1827 VSS.n420 VSS.n377 69.4405
R1828 VSS.n478 VSS.n394 69.4405
R1829 VSS.n648 VSS.n73 69.4405
R1830 VSS.n168 VSS.n152 69.4405
R1831 VSS.n178 VSS.n177 67.1161
R1832 VSS.n189 VSS.n174 67.1161
R1833 VSS.n711 VSS.n1 67.1161
R1834 VSS.n8 VSS.n6 67.1161
R1835 VSS.n703 VSS.n10 67.1161
R1836 VSS.n17 VSS.n15 67.1161
R1837 VSS.n695 VSS.n19 67.1161
R1838 VSS.n26 VSS.n24 67.1161
R1839 VSS.n687 VSS.n28 67.1161
R1840 VSS.n35 VSS.n33 67.1161
R1841 VSS.n679 VSS.n37 67.1161
R1842 VSS.n44 VSS.n42 67.1161
R1843 VSS.n671 VSS.n46 67.1161
R1844 VSS.n53 VSS.n51 67.1161
R1845 VSS.n663 VSS.n55 67.1161
R1846 VSS.n62 VSS.n60 67.1161
R1847 VSS.n555 VSS.n139 66.9639
R1848 VSS.n556 VSS.n138 66.9639
R1849 VSS.n558 VSS.n557 66.9639
R1850 VSS.n135 VSS.n134 66.9639
R1851 VSS.n564 VSS.n563 66.9639
R1852 VSS.n131 VSS.n130 66.9639
R1853 VSS.n570 VSS.n129 66.9639
R1854 VSS.n571 VSS.n128 66.9639
R1855 VSS.n574 VSS.n573 66.9639
R1856 VSS.n124 VSS.n123 66.9639
R1857 VSS.n580 VSS.n122 66.9639
R1858 VSS.n581 VSS.n121 66.9639
R1859 VSS.n584 VSS.n583 66.9639
R1860 VSS.n117 VSS.n116 66.9639
R1861 VSS.n590 VSS.n115 66.9639
R1862 VSS.n591 VSS.n114 66.9639
R1863 VSS.n594 VSS.n593 66.9639
R1864 VSS.n110 VSS.n109 66.9639
R1865 VSS.n600 VSS.n108 66.9639
R1866 VSS.n601 VSS.n107 66.9639
R1867 VSS.n604 VSS.n603 66.9639
R1868 VSS.n103 VSS.n102 66.9639
R1869 VSS.n610 VSS.n101 66.9639
R1870 VSS.n611 VSS.n100 66.9639
R1871 VSS.n614 VSS.n613 66.9639
R1872 VSS.n96 VSS.n95 66.9639
R1873 VSS.n620 VSS.n94 66.9639
R1874 VSS.n621 VSS.n93 66.9639
R1875 VSS.n624 VSS.n623 66.9639
R1876 VSS.n89 VSS.n88 66.9639
R1877 VSS.n630 VSS.n87 66.9639
R1878 VSS.n631 VSS.n86 66.9639
R1879 VSS.n634 VSS.n83 66.9639
R1880 VSS.n635 VSS.n82 66.9639
R1881 VSS.n637 VSS.n81 66.9639
R1882 VSS.n638 VSS.n80 66.9639
R1883 VSS.n165 VSS.t184 59.8776
R1884 VSS.n255 VSS.t376 59.8776
R1885 VSS.t174 VSS.n527 59.8776
R1886 VSS.n338 VSS.t46 59.8776
R1887 VSS.t233 VSS.n504 59.8776
R1888 VSS.n417 VSS.t167 59.8776
R1889 VSS.t345 VSS.n481 59.8776
R1890 VSS.t192 VSS.n651 59.8776
R1891 VSS.n170 VSS.n169 53.1823
R1892 VSS.n171 VSS.n170 53.1823
R1893 VSS.n260 VSS.n259 53.1823
R1894 VSS.n261 VSS.n260 53.1823
R1895 VSS.n523 VSS.n522 53.1823
R1896 VSS.n522 VSS.n521 53.1823
R1897 VSS.n343 VSS.n342 53.1823
R1898 VSS.n344 VSS.n343 53.1823
R1899 VSS.n500 VSS.n499 53.1823
R1900 VSS.n499 VSS.n498 53.1823
R1901 VSS.n422 VSS.n421 53.1823
R1902 VSS.n423 VSS.n422 53.1823
R1903 VSS.n477 VSS.n476 53.1823
R1904 VSS.n476 VSS.n475 53.1823
R1905 VSS.n647 VSS.n646 53.1823
R1906 VSS.n646 VSS.n645 53.1823
R1907 VSS.n167 VSS.n166 48.7505
R1908 VSS.n166 VSS.n165 48.7505
R1909 VSS.n257 VSS.n256 48.7505
R1910 VSS.n256 VSS.n255 48.7505
R1911 VSS.n526 VSS.n525 48.7505
R1912 VSS.n527 VSS.n526 48.7505
R1913 VSS.n340 VSS.n339 48.7505
R1914 VSS.n339 VSS.n338 48.7505
R1915 VSS.n503 VSS.n502 48.7505
R1916 VSS.n504 VSS.n503 48.7505
R1917 VSS.n419 VSS.n418 48.7505
R1918 VSS.n418 VSS.n417 48.7505
R1919 VSS.n480 VSS.n479 48.7505
R1920 VSS.n481 VSS.n480 48.7505
R1921 VSS.n650 VSS.n649 48.7505
R1922 VSS.n651 VSS.n650 48.7505
R1923 VSS.n252 VSS.n249 48.2672
R1924 VSS.n264 VSS.n223 48.2672
R1925 VSS.n335 VSS.n332 48.2672
R1926 VSS.n347 VSS.n306 48.2672
R1927 VSS.n414 VSS.n411 48.2672
R1928 VSS.n442 VSS.n393 48.2672
R1929 VSS.n398 VSS.n72 48.2672
R1930 VSS.n162 VSS.n159 48.2672
R1931 VSS.t40 VSS.n550 45.1409
R1932 VSS.n158 VSS.n156 45.0005
R1933 VSS.n156 VSS.n155 45.0005
R1934 VSS.n248 VSS.n245 45.0005
R1935 VSS.n245 VSS.n244 45.0005
R1936 VSS.n227 VSS.n225 45.0005
R1937 VSS.n227 VSS.n220 45.0005
R1938 VSS.n331 VSS.n328 45.0005
R1939 VSS.n328 VSS.n327 45.0005
R1940 VSS.n310 VSS.n308 45.0005
R1941 VSS.n310 VSS.n303 45.0005
R1942 VSS.n410 VSS.n407 45.0005
R1943 VSS.n407 VSS.n406 45.0005
R1944 VSS.n397 VSS.n395 45.0005
R1945 VSS.n397 VSS.n390 45.0005
R1946 VSS.n76 VSS.n74 45.0005
R1947 VSS.n76 VSS.n69 45.0005
R1948 VSS.n548 VSS.n547 39.0005
R1949 VSS.n549 VSS.n548 39.0005
R1950 VSS.n539 VSS.n538 39.0005
R1951 VSS.n540 VSS.n539 39.0005
R1952 VSS.n218 VSS.n213 39.0005
R1953 VSS.n270 VSS.n218 39.0005
R1954 VSS.n516 VSS.n515 39.0005
R1955 VSS.n517 VSS.n516 39.0005
R1956 VSS.n301 VSS.n296 39.0005
R1957 VSS.n353 VSS.n301 39.0005
R1958 VSS.n493 VSS.n492 39.0005
R1959 VSS.n494 VSS.n493 39.0005
R1960 VSS.n388 VSS.n379 39.0005
R1961 VSS.n448 VSS.n388 39.0005
R1962 VSS.n67 VSS.n66 39.0005
R1963 VSS.n404 VSS.n67 39.0005
R1964 VSS.n650 VSS.n71 34.4755
R1965 VSS.n480 VSS.n392 34.4755
R1966 VSS.n418 VSS.n409 34.4755
R1967 VSS.n503 VSS.n305 34.4755
R1968 VSS.n339 VSS.n330 34.4755
R1969 VSS.n526 VSS.n222 34.4755
R1970 VSS.n256 VSS.n247 34.4755
R1971 VSS.n166 VSS.n157 34.4755
R1972 VSS.n146 VSS.t385 31.7728
R1973 VSS.n207 VSS.t33 31.7728
R1974 VSS.n533 VSS.t60 31.7728
R1975 VSS.n290 VSS.t52 31.7728
R1976 VSS.n510 VSS.t327 31.7728
R1977 VSS.n373 VSS.t130 31.7728
R1978 VSS.n487 VSS.t142 31.7728
R1979 VSS.n384 VSS.t383 31.7728
R1980 VSS.n551 VSS.n137 28.0309
R1981 VSS.n567 VSS.n132 28.0309
R1982 VSS.n577 VSS.n125 28.0309
R1983 VSS.n587 VSS.n118 28.0309
R1984 VSS.n597 VSS.n111 28.0309
R1985 VSS.n607 VSS.n104 28.0309
R1986 VSS.n617 VSS.n97 28.0309
R1987 VSS.n627 VSS.n90 28.0309
R1988 VSS.n431 VSS.n430 28.0309
R1989 VSS.n432 VSS.n431 27.8375
R1990 VSS.n439 VSS.n90 27.8375
R1991 VSS.n426 VSS.n97 27.8375
R1992 VSS.n362 VSS.n104 27.8375
R1993 VSS.n356 VSS.n111 27.8375
R1994 VSS.n279 VSS.n118 27.8375
R1995 VSS.n273 VSS.n125 27.8375
R1996 VSS.n196 VSS.n132 27.8375
R1997 VSS.n552 VSS.n551 27.8375
R1998 VSS.n149 VSS.n148 25.9728
R1999 VSS.n150 VSS.n147 25.9728
R2000 VSS.n208 VSS.n206 25.9728
R2001 VSS.n209 VSS.n205 25.9728
R2002 VSS.n532 VSS.n214 25.9728
R2003 VSS.n531 VSS.n215 25.9728
R2004 VSS.n291 VSS.n289 25.9728
R2005 VSS.n292 VSS.n288 25.9728
R2006 VSS.n509 VSS.n297 25.9728
R2007 VSS.n508 VSS.n298 25.9728
R2008 VSS.n374 VSS.n372 25.9728
R2009 VSS.n375 VSS.n371 25.9728
R2010 VSS.n486 VSS.n380 25.9728
R2011 VSS.n485 VSS.n381 25.9728
R2012 VSS.n383 VSS.n382 25.9728
R2013 VSS.n65 VSS.n64 25.9728
R2014 VSS.n165 VSS.n155 23.1787
R2015 VSS.n255 VSS.n244 23.1787
R2016 VSS.n527 VSS.n220 23.1787
R2017 VSS.n338 VSS.n327 23.1787
R2018 VSS.n504 VSS.n303 23.1787
R2019 VSS.n417 VSS.n406 23.1787
R2020 VSS.n481 VSS.n390 23.1787
R2021 VSS.n651 VSS.n69 23.1787
R2022 VSS.n249 VSS.n203 23.1494
R2023 VSS.n267 VSS.n223 23.1494
R2024 VSS.n332 VSS.n286 23.1494
R2025 VSS.n350 VSS.n306 23.1494
R2026 VSS.n411 VSS.n369 23.1494
R2027 VSS.n445 VSS.n393 23.1494
R2028 VSS.n401 VSS.n72 23.1494
R2029 VSS.n159 VSS.n145 23.1494
R2030 VSS.n545 VSS.n544 22.5005
R2031 VSS.n544 VSS.n543 22.5005
R2032 VSS.n536 VSS.n212 22.5005
R2033 VSS.n262 VSS.n212 22.5005
R2034 VSS.n219 VSS.n217 22.5005
R2035 VSS.n520 VSS.n219 22.5005
R2036 VSS.n513 VSS.n295 22.5005
R2037 VSS.n345 VSS.n295 22.5005
R2038 VSS.n302 VSS.n300 22.5005
R2039 VSS.n497 VSS.n302 22.5005
R2040 VSS.n490 VSS.n378 22.5005
R2041 VSS.n424 VSS.n378 22.5005
R2042 VSS.n389 VSS.n387 22.5005
R2043 VSS.n474 VSS.n389 22.5005
R2044 VSS.n68 VSS.n63 22.5005
R2045 VSS.n644 VSS.n68 22.5005
R2046 VSS.n464 VSS.n461 19.761
R2047 VSS.n456 VSS.n453 19.761
R2048 VSS.n316 VSS.n315 19.761
R2049 VSS.n324 VSS.n321 19.761
R2050 VSS.n233 VSS.n232 19.761
R2051 VSS.n241 VSS.n238 19.761
R2052 VSS.n183 VSS.n182 19.761
R2053 VSS.n469 VSS.n468 19.761
R2054 VSS.n536 VSS.n211 18.2672
R2055 VSS.n224 VSS.n217 18.2672
R2056 VSS.n513 VSS.n294 18.2672
R2057 VSS.n307 VSS.n300 18.2672
R2058 VSS.n490 VSS.n377 18.2672
R2059 VSS.n394 VSS.n387 18.2672
R2060 VSS.n73 VSS.n63 18.2672
R2061 VSS.n545 VSS.n152 18.2672
R2062 VSS.n177 VSS.t263 17.4005
R2063 VSS.n177 VSS.t261 17.4005
R2064 VSS.n174 VSS.t331 17.4005
R2065 VSS.n174 VSS.t304 17.4005
R2066 VSS.n1 VSS.t325 17.4005
R2067 VSS.n1 VSS.t15 17.4005
R2068 VSS.n6 VSS.t235 17.4005
R2069 VSS.n6 VSS.t297 17.4005
R2070 VSS.n10 VSS.t339 17.4005
R2071 VSS.n10 VSS.t281 17.4005
R2072 VSS.n15 VSS.t187 17.4005
R2073 VSS.n15 VSS.t202 17.4005
R2074 VSS.n19 VSS.t64 17.4005
R2075 VSS.n19 VSS.t153 17.4005
R2076 VSS.n24 VSS.t17 17.4005
R2077 VSS.n24 VSS.t177 17.4005
R2078 VSS.n28 VSS.t210 17.4005
R2079 VSS.n28 VSS.t212 17.4005
R2080 VSS.n33 VSS.t189 17.4005
R2081 VSS.n33 VSS.t285 17.4005
R2082 VSS.n37 VSS.t62 17.4005
R2083 VSS.n37 VSS.t191 17.4005
R2084 VSS.n42 VSS.t289 17.4005
R2085 VSS.n42 VSS.t250 17.4005
R2086 VSS.n46 VSS.t258 17.4005
R2087 VSS.n46 VSS.t91 17.4005
R2088 VSS.n51 VSS.t79 17.4005
R2089 VSS.n51 VSS.t227 17.4005
R2090 VSS.n55 VSS.t31 17.4005
R2091 VSS.n55 VSS.t69 17.4005
R2092 VSS.n60 VSS.t71 17.4005
R2093 VSS.n60 VSS.t344 17.4005
R2094 VSS.n139 VSS.t266 17.4005
R2095 VSS.n139 VSS.t155 17.4005
R2096 VSS.n138 VSS.t283 17.4005
R2097 VSS.n138 VSS.t77 17.4005
R2098 VSS.n557 VSS.t380 17.4005
R2099 VSS.n557 VSS.t29 17.4005
R2100 VSS.n134 VSS.t273 17.4005
R2101 VSS.n134 VSS.t41 17.4005
R2102 VSS.n563 VSS.t389 17.4005
R2103 VSS.n563 VSS.t223 17.4005
R2104 VSS.n130 VSS.t352 17.4005
R2105 VSS.n130 VSS.t25 17.4005
R2106 VSS.n129 VSS.t160 17.4005
R2107 VSS.n129 VSS.t378 17.4005
R2108 VSS.n128 VSS.t214 17.4005
R2109 VSS.n128 VSS.t81 17.4005
R2110 VSS.n573 VSS.t9 17.4005
R2111 VSS.n573 VSS.t337 17.4005
R2112 VSS.n123 VSS.t95 17.4005
R2113 VSS.n123 VSS.t147 17.4005
R2114 VSS.n122 VSS.t157 17.4005
R2115 VSS.n122 VSS.t27 17.4005
R2116 VSS.n121 VSS.t347 17.4005
R2117 VSS.n121 VSS.t48 17.4005
R2118 VSS.n583 VSS.t268 17.4005
R2119 VSS.n583 VSS.t45 17.4005
R2120 VSS.n116 VSS.t246 17.4005
R2121 VSS.n116 VSS.t373 17.4005
R2122 VSS.n115 VSS.t232 17.4005
R2123 VSS.n115 VSS.t230 17.4005
R2124 VSS.n114 VSS.t200 17.4005
R2125 VSS.n114 VSS.t240 17.4005
R2126 VSS.n593 VSS.t144 17.4005
R2127 VSS.n593 VSS.t391 17.4005
R2128 VSS.n109 VSS.t208 17.4005
R2129 VSS.n109 VSS.t287 17.4005
R2130 VSS.n108 VSS.t329 17.4005
R2131 VSS.n108 VSS.t98 17.4005
R2132 VSS.n107 VSS.t369 17.4005
R2133 VSS.n107 VSS.t366 17.4005
R2134 VSS.n603 VSS.t248 17.4005
R2135 VSS.n603 VSS.t164 17.4005
R2136 VSS.n102 VSS.t238 17.4005
R2137 VSS.n102 VSS.t350 17.4005
R2138 VSS.n101 VSS.t116 17.4005
R2139 VSS.n101 VSS.t295 17.4005
R2140 VSS.n100 VSS.t399 17.4005
R2141 VSS.n100 VSS.t395 17.4005
R2142 VSS.n613 VSS.t124 17.4005
R2143 VSS.n613 VSS.t120 17.4005
R2144 VSS.n95 VSS.t126 17.4005
R2145 VSS.n95 VSS.t122 17.4005
R2146 VSS.n94 VSS.t3 17.4005
R2147 VSS.n94 VSS.t6 17.4005
R2148 VSS.n93 VSS.t19 17.4005
R2149 VSS.n93 VSS.t1 17.4005
R2150 VSS.n623 VSS.t108 17.4005
R2151 VSS.n623 VSS.t111 17.4005
R2152 VSS.n88 VSS.t105 17.4005
R2153 VSS.n88 VSS.t113 17.4005
R2154 VSS.n87 VSS.t319 17.4005
R2155 VSS.n87 VSS.t321 17.4005
R2156 VSS.n86 VSS.t252 17.4005
R2157 VSS.n86 VSS.t316 17.4005
R2158 VSS.n83 VSS.t314 17.4005
R2159 VSS.n83 VSS.t310 17.4005
R2160 VSS.n82 VSS.t312 17.4005
R2161 VSS.n82 VSS.t308 17.4005
R2162 VSS.n81 VSS.t172 17.4005
R2163 VSS.n81 VSS.t293 17.4005
R2164 VSS.n80 VSS.t302 17.4005
R2165 VSS.n80 VSS.t291 17.4005
R2166 VSS.n668 VSS.n48 17.2064
R2167 VSS.n461 VSS.n48 17.2064
R2168 VSS.n676 VSS.n39 17.2064
R2169 VSS.n453 VSS.n39 17.2064
R2170 VSS.n684 VSS.n30 17.2064
R2171 VSS.n316 VSS.n30 17.2064
R2172 VSS.n692 VSS.n21 17.2064
R2173 VSS.n321 VSS.n21 17.2064
R2174 VSS.n700 VSS.n12 17.2064
R2175 VSS.n233 VSS.n12 17.2064
R2176 VSS.n708 VSS.n3 17.2064
R2177 VSS.n238 VSS.n3 17.2064
R2178 VSS.n185 VSS.n184 17.2064
R2179 VSS.n184 VSS.n183 17.2064
R2180 VSS.n660 VSS.n57 17.2064
R2181 VSS.n469 VSS.n57 17.2064
R2182 VSS.n546 VSS.n144 15.3952
R2183 VSS.t93 VSS.n144 15.3952
R2184 VSS.n537 VSS.n202 15.3952
R2185 VSS.t128 VSS.n202 15.3952
R2186 VSS.n529 VSS.n528 15.3952
R2187 VSS.n528 VSS.t10 15.3952
R2188 VSS.n514 VSS.n285 15.3952
R2189 VSS.t179 VSS.n285 15.3952
R2190 VSS.n506 VSS.n505 15.3952
R2191 VSS.n505 VSS.t175 15.3952
R2192 VSS.n491 VSS.n368 15.3952
R2193 VSS.t162 VSS.n368 15.3952
R2194 VSS.n483 VSS.n482 15.3952
R2195 VSS.n482 VSS.t7 15.3952
R2196 VSS.n653 VSS.n652 15.3952
R2197 VSS.n652 VSS.t42 15.3952
R2198 VSS VSS.n656 6.94083
R2199 VSS.n148 VSS.t54 5.8005
R2200 VSS.n148 VSS.t362 5.8005
R2201 VSS.n147 VSS.t358 5.8005
R2202 VSS.n147 VSS.t393 5.8005
R2203 VSS.n206 VSS.t256 5.8005
R2204 VSS.n206 VSS.t56 5.8005
R2205 VSS.n205 VSS.t364 5.8005
R2206 VSS.n205 VSS.t360 5.8005
R2207 VSS.n214 VSS.t35 5.8005
R2208 VSS.n214 VSS.t140 5.8005
R2209 VSS.n215 VSS.t89 5.8005
R2210 VSS.n215 VSS.t387 5.8005
R2211 VSS.n289 VSS.t216 5.8005
R2212 VSS.n289 VSS.t136 5.8005
R2213 VSS.n288 VSS.t244 5.8005
R2214 VSS.n288 VSS.t50 5.8005
R2215 VSS.n297 VSS.t218 5.8005
R2216 VSS.n297 VSS.t138 5.8005
R2217 VSS.n298 VSS.t342 5.8005
R2218 VSS.n298 VSS.t58 5.8005
R2219 VSS.n372 VSS.t242 5.8005
R2220 VSS.n372 VSS.t87 5.8005
R2221 VSS.n371 VSS.t83 5.8005
R2222 VSS.n371 VSS.t220 5.8005
R2223 VSS.n380 VSS.t149 5.8005
R2224 VSS.n380 VSS.t37 5.8005
R2225 VSS.n381 VSS.t254 5.8005
R2226 VSS.n381 VSS.t85 5.8005
R2227 VSS.n382 VSS.t13 5.8005
R2228 VSS.n382 VSS.t183 5.8005
R2229 VSS.n64 VSS.t39 5.8005
R2230 VSS.n64 VSS.t275 5.8005
R2231 VSS.n184 VSS.n172 5.79462
R2232 VSS.n239 VSS.n3 5.79462
R2233 VSS.n230 VSS.n12 5.79462
R2234 VSS.n322 VSS.n21 5.79462
R2235 VSS.n313 VSS.n30 5.79462
R2236 VSS.n454 VSS.n39 5.79462
R2237 VSS.n462 VSS.n48 5.79462
R2238 VSS.n466 VSS.n57 5.79462
R2239 VSS.n656 VSS 4.62996
R2240 VSS.n656 VSS 4.34685
R2241 VSS.n171 VSS.n155 3.86354
R2242 VSS.n261 VSS.n244 3.86354
R2243 VSS.n521 VSS.n220 3.86354
R2244 VSS.n344 VSS.n327 3.86354
R2245 VSS.n498 VSS.n303 3.86354
R2246 VSS.n423 VSS.n406 3.86354
R2247 VSS.n475 VSS.n390 3.86354
R2248 VSS.n645 VSS.n69 3.86354
R2249 VSS.n555 VSS.n554 3.0429
R2250 VSS.n551 VSS.n140 2.96352
R2251 VSS.n197 VSS.n132 2.96352
R2252 VSS.n274 VSS.n125 2.96352
R2253 VSS.n280 VSS.n118 2.96352
R2254 VSS.n357 VSS.n111 2.96352
R2255 VSS.n363 VSS.n104 2.96352
R2256 VSS.n427 VSS.n97 2.96352
R2257 VSS.n436 VSS.n90 2.96352
R2258 VSS.n431 VSS.n78 2.96352
R2259 VSS.n566 VSS.n565 2.7955
R2260 VSS.n572 VSS.n127 2.7955
R2261 VSS.n576 VSS.n575 2.7955
R2262 VSS.n582 VSS.n120 2.7955
R2263 VSS.n586 VSS.n585 2.7955
R2264 VSS.n592 VSS.n113 2.7955
R2265 VSS.n596 VSS.n595 2.7955
R2266 VSS.n602 VSS.n106 2.7955
R2267 VSS.n606 VSS.n605 2.7955
R2268 VSS.n612 VSS.n99 2.7955
R2269 VSS.n616 VSS.n615 2.7955
R2270 VSS.n622 VSS.n92 2.7955
R2271 VSS.n626 VSS.n625 2.7955
R2272 VSS.n632 VSS.n85 2.7955
R2273 VSS.n633 VSS.n84 2.7955
R2274 VSS.n640 VSS.n639 2.7955
R2275 VSS.n562 VSS.n561 2.7955
R2276 VSS.n179 VSS.n178 2.60207
R2277 VSS.n187 VSS.n175 2.39175
R2278 VSS.n4 VSS.n2 2.39175
R2279 VSS.n13 VSS.n11 2.39175
R2280 VSS.n22 VSS.n20 2.39175
R2281 VSS.n31 VSS.n29 2.39175
R2282 VSS.n40 VSS.n38 2.39175
R2283 VSS.n49 VSS.n47 2.39175
R2284 VSS.n58 VSS.n56 2.39175
R2285 VSS.n191 VSS.n190 2.3631
R2286 VSS.n712 VSS.n0 2.3631
R2287 VSS.n706 VSS.n705 2.3631
R2288 VSS.n704 VSS.n9 2.3631
R2289 VSS.n698 VSS.n697 2.3631
R2290 VSS.n696 VSS.n18 2.3631
R2291 VSS.n690 VSS.n689 2.3631
R2292 VSS.n688 VSS.n27 2.3631
R2293 VSS.n682 VSS.n681 2.3631
R2294 VSS.n680 VSS.n36 2.3631
R2295 VSS.n674 VSS.n673 2.3631
R2296 VSS.n672 VSS.n45 2.3631
R2297 VSS.n666 VSS.n665 2.3631
R2298 VSS.n664 VSS.n54 2.3631
R2299 VSS.n658 VSS.n657 2.3631
R2300 VSS.n258 VSS.n257 2.2405
R2301 VSS.n525 VSS.n524 2.2405
R2302 VSS.n341 VSS.n340 2.2405
R2303 VSS.n502 VSS.n501 2.2405
R2304 VSS.n420 VSS.n419 2.2405
R2305 VSS.n479 VSS.n478 2.2405
R2306 VSS.n649 VSS.n648 2.2405
R2307 VSS.n168 VSS.n167 2.2405
R2308 VSS.t357 VSS.n164 1.93202
R2309 VSS.t363 VSS.n254 1.93202
R2310 VSS.n266 VSS.t88 1.93202
R2311 VSS.t243 VSS.n337 1.93202
R2312 VSS.n349 VSS.t341 1.93202
R2313 VSS.t82 VSS.n416 1.93202
R2314 VSS.n444 VSS.t253 1.93202
R2315 VSS.n400 VSS.t38 1.93202
R2316 VSS.n545 VSS.n153 1.56378
R2317 VSS.n536 VSS.n535 1.56378
R2318 VSS.n217 VSS.n216 1.56378
R2319 VSS.n513 VSS.n512 1.56378
R2320 VSS.n300 VSS.n299 1.56378
R2321 VSS.n490 VSS.n489 1.56378
R2322 VSS.n387 VSS.n386 1.56378
R2323 VSS.n655 VSS.n63 1.56378
R2324 VSS.n547 VSS.n146 1.51802
R2325 VSS.n565 VSS 1.3768
R2326 VSS.n575 VSS 1.3768
R2327 VSS.n585 VSS 1.3768
R2328 VSS.n595 VSS 1.3768
R2329 VSS.n605 VSS 1.3768
R2330 VSS.n615 VSS 1.3768
R2331 VSS.n625 VSS 1.3768
R2332 VSS.n633 VSS 1.3768
R2333 VSS.n538 VSS.n204 1.37182
R2334 VSS.n534 VSS.n213 1.37182
R2335 VSS.n515 VSS.n287 1.37182
R2336 VSS.n511 VSS.n296 1.37182
R2337 VSS.n492 VSS.n370 1.37182
R2338 VSS.n488 VSS.n379 1.37182
R2339 VSS.n385 VSS.n66 1.37182
R2340 VSS.n568 VSS.n567 0.8005
R2341 VSS.n578 VSS.n577 0.8005
R2342 VSS.n588 VSS.n587 0.8005
R2343 VSS.n598 VSS.n597 0.8005
R2344 VSS.n608 VSS.n607 0.8005
R2345 VSS.n618 VSS.n617 0.8005
R2346 VSS.n628 VSS.n627 0.8005
R2347 VSS.n430 VSS.n79 0.8005
R2348 VSS.n560 VSS.n137 0.8005
R2349 VSS.n153 VSS.n151 0.785098
R2350 VSS.n535 VSS.n210 0.785098
R2351 VSS.n530 VSS.n216 0.785098
R2352 VSS.n512 VSS.n293 0.785098
R2353 VSS.n507 VSS.n299 0.785098
R2354 VSS.n489 VSS.n376 0.785098
R2355 VSS.n484 VSS.n386 0.785098
R2356 VSS.n655 VSS.n654 0.785098
R2357 VSS VSS.n712 0.669618
R2358 VSS VSS.n704 0.669618
R2359 VSS VSS.n696 0.669618
R2360 VSS VSS.n688 0.669618
R2361 VSS VSS.n680 0.669618
R2362 VSS VSS.n672 0.669618
R2363 VSS VSS.n664 0.669618
R2364 VSS.n186 VSS.n185 0.58175
R2365 VSS.n709 VSS.n708 0.58175
R2366 VSS.n701 VSS.n700 0.58175
R2367 VSS.n693 VSS.n692 0.58175
R2368 VSS.n685 VSS.n684 0.58175
R2369 VSS.n677 VSS.n676 0.58175
R2370 VSS.n669 VSS.n668 0.58175
R2371 VSS.n661 VSS.n660 0.58175
R2372 VSS.n569 VSS.n568 0.547559
R2373 VSS.n579 VSS.n578 0.547559
R2374 VSS.n589 VSS.n588 0.547559
R2375 VSS.n599 VSS.n598 0.547559
R2376 VSS.n609 VSS.n608 0.547559
R2377 VSS.n619 VSS.n618 0.547559
R2378 VSS.n629 VSS.n628 0.547559
R2379 VSS.n636 VSS.n79 0.547559
R2380 VSS.n560 VSS.n559 0.547559
R2381 VSS VSS.n153 0.522821
R2382 VSS.n535 VSS 0.522821
R2383 VSS VSS.n216 0.522821
R2384 VSS.n512 VSS 0.522821
R2385 VSS VSS.n299 0.522821
R2386 VSS.n489 VSS 0.522821
R2387 VSS.n386 VSS 0.522821
R2388 VSS VSS.n655 0.522821
R2389 VSS.n537 VSS.n210 0.517167
R2390 VSS.n530 VSS.n529 0.517167
R2391 VSS.n514 VSS.n293 0.517167
R2392 VSS.n507 VSS.n506 0.517167
R2393 VSS.n491 VSS.n376 0.517167
R2394 VSS.n484 VSS.n483 0.517167
R2395 VSS.n654 VSS.n653 0.517167
R2396 VSS.n546 VSS.n151 0.517167
R2397 VSS.n204 VSS 0.455857
R2398 VSS VSS.n534 0.455857
R2399 VSS.n287 VSS 0.455857
R2400 VSS VSS.n511 0.455857
R2401 VSS.n370 VSS 0.455857
R2402 VSS VSS.n488 0.455857
R2403 VSS VSS.n385 0.455857
R2404 VSS.n185 VSS.n173 0.376971
R2405 VSS.n708 VSS.n707 0.376971
R2406 VSS.n700 VSS.n699 0.376971
R2407 VSS.n692 VSS.n691 0.376971
R2408 VSS.n684 VSS.n683 0.376971
R2409 VSS.n676 VSS.n675 0.376971
R2410 VSS.n668 VSS.n667 0.376971
R2411 VSS.n660 VSS.n659 0.376971
R2412 VSS.n178 VSS.n176 0.324029
R2413 VSS.n189 VSS.n188 0.324029
R2414 VSS.n711 VSS.n710 0.324029
R2415 VSS.n8 VSS.n7 0.324029
R2416 VSS.n703 VSS.n702 0.324029
R2417 VSS.n17 VSS.n16 0.324029
R2418 VSS.n695 VSS.n694 0.324029
R2419 VSS.n26 VSS.n25 0.324029
R2420 VSS.n687 VSS.n686 0.324029
R2421 VSS.n35 VSS.n34 0.324029
R2422 VSS.n679 VSS.n678 0.324029
R2423 VSS.n44 VSS.n43 0.324029
R2424 VSS.n671 VSS.n670 0.324029
R2425 VSS.n53 VSS.n52 0.324029
R2426 VSS.n663 VSS.n662 0.324029
R2427 VSS.n62 VSS.n61 0.324029
R2428 VSS.n559 VSS.n556 0.255708
R2429 VSS.n569 VSS.n131 0.255708
R2430 VSS.n579 VSS.n124 0.255708
R2431 VSS.n589 VSS.n117 0.255708
R2432 VSS.n599 VSS.n110 0.255708
R2433 VSS.n609 VSS.n103 0.255708
R2434 VSS.n619 VSS.n96 0.255708
R2435 VSS.n629 VSS.n89 0.255708
R2436 VSS.n636 VSS.n635 0.255708
R2437 VSS.n562 VSS.n135 0.247896
R2438 VSS.n565 VSS.n564 0.247896
R2439 VSS.n572 VSS.n571 0.247896
R2440 VSS.n575 VSS.n574 0.247896
R2441 VSS.n582 VSS.n581 0.247896
R2442 VSS.n585 VSS.n584 0.247896
R2443 VSS.n592 VSS.n591 0.247896
R2444 VSS.n595 VSS.n594 0.247896
R2445 VSS.n602 VSS.n601 0.247896
R2446 VSS.n605 VSS.n604 0.247896
R2447 VSS.n612 VSS.n611 0.247896
R2448 VSS.n615 VSS.n614 0.247896
R2449 VSS.n622 VSS.n621 0.247896
R2450 VSS.n625 VSS.n624 0.247896
R2451 VSS.n632 VSS.n631 0.247896
R2452 VSS.n634 VSS.n633 0.247896
R2453 VSS.n639 VSS.n638 0.247896
R2454 VSS.n151 VSS.n150 0.246036
R2455 VSS.n210 VSS.n209 0.246036
R2456 VSS.n531 VSS.n530 0.246036
R2457 VSS.n293 VSS.n292 0.246036
R2458 VSS.n508 VSS.n507 0.246036
R2459 VSS.n376 VSS.n375 0.246036
R2460 VSS.n485 VSS.n484 0.246036
R2461 VSS.n654 VSS.n65 0.246036
R2462 VSS.n559 VSS.n558 0.240083
R2463 VSS.n570 VSS.n569 0.240083
R2464 VSS.n580 VSS.n579 0.240083
R2465 VSS.n590 VSS.n589 0.240083
R2466 VSS.n600 VSS.n599 0.240083
R2467 VSS.n610 VSS.n609 0.240083
R2468 VSS.n620 VSS.n619 0.240083
R2469 VSS.n630 VSS.n629 0.240083
R2470 VSS.n637 VSS.n636 0.240083
R2471 VSS.n712 VSS.n711 0.239471
R2472 VSS.n704 VSS.n703 0.239471
R2473 VSS.n696 VSS.n695 0.239471
R2474 VSS.n688 VSS.n687 0.239471
R2475 VSS.n680 VSS.n679 0.239471
R2476 VSS.n672 VSS.n671 0.239471
R2477 VSS.n664 VSS.n663 0.239471
R2478 VSS.n190 VSS.n189 0.232118
R2479 VSS.n705 VSS.n8 0.232118
R2480 VSS.n697 VSS.n17 0.232118
R2481 VSS.n689 VSS.n26 0.232118
R2482 VSS.n681 VSS.n35 0.232118
R2483 VSS.n673 VSS.n44 0.232118
R2484 VSS.n665 VSS.n53 0.232118
R2485 VSS.n657 VSS.n62 0.232118
R2486 VSS.n556 VSS.n555 0.229667
R2487 VSS.n558 VSS.n135 0.229667
R2488 VSS.n564 VSS.n131 0.229667
R2489 VSS.n571 VSS.n570 0.229667
R2490 VSS.n574 VSS.n124 0.229667
R2491 VSS.n581 VSS.n580 0.229667
R2492 VSS.n584 VSS.n117 0.229667
R2493 VSS.n591 VSS.n590 0.229667
R2494 VSS.n594 VSS.n110 0.229667
R2495 VSS.n601 VSS.n600 0.229667
R2496 VSS.n604 VSS.n103 0.229667
R2497 VSS.n611 VSS.n610 0.229667
R2498 VSS.n614 VSS.n96 0.229667
R2499 VSS.n621 VSS.n620 0.229667
R2500 VSS.n624 VSS.n89 0.229667
R2501 VSS.n631 VSS.n630 0.229667
R2502 VSS.n635 VSS.n634 0.229667
R2503 VSS.n638 VSS.n637 0.229667
R2504 VSS.n149 VSS.n146 0.196929
R2505 VSS.n150 VSS.n149 0.196929
R2506 VSS.n208 VSS.n207 0.196929
R2507 VSS.n209 VSS.n208 0.196929
R2508 VSS.n533 VSS.n532 0.196929
R2509 VSS.n532 VSS.n531 0.196929
R2510 VSS.n291 VSS.n290 0.196929
R2511 VSS.n292 VSS.n291 0.196929
R2512 VSS.n510 VSS.n509 0.196929
R2513 VSS.n509 VSS.n508 0.196929
R2514 VSS.n374 VSS.n373 0.196929
R2515 VSS.n375 VSS.n374 0.196929
R2516 VSS.n487 VSS.n486 0.196929
R2517 VSS.n486 VSS.n485 0.196929
R2518 VSS.n384 VSS.n383 0.196929
R2519 VSS.n383 VSS.n65 0.196929
R2520 VSS VSS.n562 0.147635
R2521 VSS VSS.n572 0.147635
R2522 VSS VSS.n582 0.147635
R2523 VSS VSS.n592 0.147635
R2524 VSS VSS.n602 0.147635
R2525 VSS VSS.n612 0.147635
R2526 VSS VSS.n622 0.147635
R2527 VSS VSS.n632 0.147635
R2528 VSS.n639 VSS 0.147635
R2529 VSS.n207 VSS.n204 0.146705
R2530 VSS.n534 VSS.n533 0.146705
R2531 VSS.n290 VSS.n287 0.146705
R2532 VSS.n511 VSS.n510 0.146705
R2533 VSS.n373 VSS.n370 0.146705
R2534 VSS.n488 VSS.n487 0.146705
R2535 VSS.n385 VSS.n384 0.146705
R2536 VSS.n188 VSS.n187 0.124275
R2537 VSS.n7 VSS.n2 0.124275
R2538 VSS.n16 VSS.n11 0.124275
R2539 VSS.n25 VSS.n20 0.124275
R2540 VSS.n34 VSS.n29 0.124275
R2541 VSS.n43 VSS.n38 0.124275
R2542 VSS.n52 VSS.n47 0.124275
R2543 VSS.n61 VSS.n56 0.124275
R2544 VSS.n186 VSS.n176 0.120598
R2545 VSS.n710 VSS.n709 0.120598
R2546 VSS.n702 VSS.n701 0.120598
R2547 VSS.n694 VSS.n693 0.120598
R2548 VSS.n686 VSS.n685 0.120598
R2549 VSS.n678 VSS.n677 0.120598
R2550 VSS.n670 VSS.n669 0.120598
R2551 VSS.n662 VSS.n661 0.120598
R2552 VSS.n190 VSS 0.113245
R2553 VSS.n705 VSS 0.113245
R2554 VSS.n697 VSS 0.113245
R2555 VSS.n689 VSS 0.113245
R2556 VSS.n681 VSS 0.113245
R2557 VSS.n673 VSS 0.113245
R2558 VSS.n665 VSS 0.113245
R2559 VSS.n657 VSS 0.113245
R2560 VSS.n187 VSS.n186 0.00417647
R2561 VSS.n709 VSS.n2 0.00417647
R2562 VSS.n701 VSS.n11 0.00417647
R2563 VSS.n693 VSS.n20 0.00417647
R2564 VSS.n685 VSS.n29 0.00417647
R2565 VSS.n677 VSS.n38 0.00417647
R2566 VSS.n669 VSS.n47 0.00417647
R2567 VSS.n661 VSS.n56 0.00417647
R2568 stop_strong.n0 stop_strong.t25 851.506
R2569 stop_strong.n6 stop_strong.t15 851.506
R2570 stop_strong.n13 stop_strong.t49 851.506
R2571 stop_strong.n20 stop_strong.t28 851.506
R2572 stop_strong.n27 stop_strong.t19 851.506
R2573 stop_strong.n34 stop_strong.t6 851.506
R2574 stop_strong.n41 stop_strong.t22 851.506
R2575 stop_strong.n48 stop_strong.t18 851.506
R2576 stop_strong.n0 stop_strong.t27 850.414
R2577 stop_strong.n6 stop_strong.t55 850.414
R2578 stop_strong.n13 stop_strong.t45 850.414
R2579 stop_strong.n20 stop_strong.t34 850.414
R2580 stop_strong.n27 stop_strong.t35 850.414
R2581 stop_strong.n34 stop_strong.t31 850.414
R2582 stop_strong.n41 stop_strong.t23 850.414
R2583 stop_strong.n48 stop_strong.t13 850.414
R2584 stop_strong.n1 stop_strong.t44 665.16
R2585 stop_strong.n7 stop_strong.t33 665.16
R2586 stop_strong.n14 stop_strong.t3 665.16
R2587 stop_strong.n21 stop_strong.t52 665.16
R2588 stop_strong.n28 stop_strong.t38 665.16
R2589 stop_strong.n35 stop_strong.t7 665.16
R2590 stop_strong.n42 stop_strong.t41 665.16
R2591 stop_strong.n49 stop_strong.t30 665.16
R2592 stop_strong.n1 stop_strong.t32 523.774
R2593 stop_strong.n2 stop_strong.t8 523.774
R2594 stop_strong.n3 stop_strong.t42 523.774
R2595 stop_strong.n4 stop_strong.t2 523.774
R2596 stop_strong.n7 stop_strong.t9 523.774
R2597 stop_strong.n8 stop_strong.t43 523.774
R2598 stop_strong.n9 stop_strong.t17 523.774
R2599 stop_strong.n10 stop_strong.t50 523.774
R2600 stop_strong.n14 stop_strong.t37 523.774
R2601 stop_strong.n15 stop_strong.t0 523.774
R2602 stop_strong.n16 stop_strong.t51 523.774
R2603 stop_strong.n17 stop_strong.t39 523.774
R2604 stop_strong.n21 stop_strong.t11 523.774
R2605 stop_strong.n22 stop_strong.t46 523.774
R2606 stop_strong.n23 stop_strong.t20 523.774
R2607 stop_strong.n24 stop_strong.t53 523.774
R2608 stop_strong.n28 stop_strong.t12 523.774
R2609 stop_strong.n29 stop_strong.t47 523.774
R2610 stop_strong.n30 stop_strong.t21 523.774
R2611 stop_strong.n31 stop_strong.t54 523.774
R2612 stop_strong.n35 stop_strong.t40 523.774
R2613 stop_strong.n36 stop_strong.t36 523.774
R2614 stop_strong.n37 stop_strong.t10 523.774
R2615 stop_strong.n38 stop_strong.t29 523.774
R2616 stop_strong.n42 stop_strong.t16 523.774
R2617 stop_strong.n43 stop_strong.t4 523.774
R2618 stop_strong.n44 stop_strong.t24 523.774
R2619 stop_strong.n45 stop_strong.t1 523.774
R2620 stop_strong.n49 stop_strong.t5 523.774
R2621 stop_strong.n50 stop_strong.t26 523.774
R2622 stop_strong.n51 stop_strong.t14 523.774
R2623 stop_strong.n52 stop_strong.t48 523.774
R2624 stop_strong.n5 stop_strong.n4 213.51
R2625 stop_strong.n11 stop_strong.n10 213.51
R2626 stop_strong.n18 stop_strong.n17 213.51
R2627 stop_strong.n25 stop_strong.n24 213.51
R2628 stop_strong.n32 stop_strong.n31 213.51
R2629 stop_strong.n39 stop_strong.n38 213.51
R2630 stop_strong.n46 stop_strong.n45 213.51
R2631 stop_strong.n53 stop_strong.n52 213.51
R2632 stop_strong.n4 stop_strong.n3 141.387
R2633 stop_strong.n3 stop_strong.n2 141.387
R2634 stop_strong.n2 stop_strong.n1 141.387
R2635 stop_strong.n10 stop_strong.n9 141.387
R2636 stop_strong.n9 stop_strong.n8 141.387
R2637 stop_strong.n8 stop_strong.n7 141.387
R2638 stop_strong.n17 stop_strong.n16 141.387
R2639 stop_strong.n16 stop_strong.n15 141.387
R2640 stop_strong.n15 stop_strong.n14 141.387
R2641 stop_strong.n24 stop_strong.n23 141.387
R2642 stop_strong.n23 stop_strong.n22 141.387
R2643 stop_strong.n22 stop_strong.n21 141.387
R2644 stop_strong.n31 stop_strong.n30 141.387
R2645 stop_strong.n30 stop_strong.n29 141.387
R2646 stop_strong.n29 stop_strong.n28 141.387
R2647 stop_strong.n38 stop_strong.n37 141.387
R2648 stop_strong.n37 stop_strong.n36 141.387
R2649 stop_strong.n36 stop_strong.n35 141.387
R2650 stop_strong.n45 stop_strong.n44 141.387
R2651 stop_strong.n44 stop_strong.n43 141.387
R2652 stop_strong.n43 stop_strong.n42 141.387
R2653 stop_strong.n52 stop_strong.n51 141.387
R2654 stop_strong.n51 stop_strong.n50 141.387
R2655 stop_strong.n50 stop_strong.n49 141.387
R2656 stop_strong stop_strong.n5 11.8482
R2657 stop_strong.n12 stop_strong.n11 9.66066
R2658 stop_strong.n19 stop_strong.n18 9.66066
R2659 stop_strong.n26 stop_strong.n25 9.66066
R2660 stop_strong.n33 stop_strong.n32 9.66066
R2661 stop_strong.n40 stop_strong.n39 9.66066
R2662 stop_strong.n47 stop_strong.n46 9.66066
R2663 stop_strong.n54 stop_strong.n53 9.66066
R2664 stop_strong stop_strong.n12 2.188
R2665 stop_strong stop_strong.n19 2.188
R2666 stop_strong stop_strong.n26 2.188
R2667 stop_strong stop_strong.n33 2.188
R2668 stop_strong stop_strong.n40 2.188
R2669 stop_strong stop_strong.n47 2.188
R2670 stop_strong.n54 stop_strong 2.188
R2671 stop_strong.n5 stop_strong.n0 1.05649
R2672 stop_strong.n11 stop_strong.n6 1.05649
R2673 stop_strong.n18 stop_strong.n13 1.05649
R2674 stop_strong.n25 stop_strong.n20 1.05649
R2675 stop_strong.n32 stop_strong.n27 1.05649
R2676 stop_strong.n39 stop_strong.n34 1.05649
R2677 stop_strong.n46 stop_strong.n41 1.05649
R2678 stop_strong.n53 stop_strong.n48 1.05649
R2679 stop_strong.n12 stop_strong 0.6655
R2680 stop_strong.n19 stop_strong 0.6655
R2681 stop_strong.n26 stop_strong 0.6655
R2682 stop_strong.n33 stop_strong 0.6655
R2683 stop_strong.n40 stop_strong 0.6655
R2684 stop_strong.n47 stop_strong 0.6655
R2685 stop_strong stop_strong.n54 0.6655
R2686 a_11980_2192.n4 a_11980_2192.t0 32.0282
R2687 a_11980_2192.n9 a_11980_2192.n0 25.7663
R2688 a_11980_2192.n6 a_11980_2192.n1 25.75
R2689 a_11980_2192.n5 a_11980_2192.n2 25.75
R2690 a_11980_2192.n4 a_11980_2192.n3 25.75
R2691 a_11980_2192.n10 a_11980_2192.n9 25.288
R2692 a_11980_2192.n8 a_11980_2192.n7 24.288
R2693 a_11980_2192.n7 a_11980_2192.t9 5.8005
R2694 a_11980_2192.n7 a_11980_2192.t11 5.8005
R2695 a_11980_2192.n1 a_11980_2192.t12 5.8005
R2696 a_11980_2192.n1 a_11980_2192.t5 5.8005
R2697 a_11980_2192.n2 a_11980_2192.t4 5.8005
R2698 a_11980_2192.n2 a_11980_2192.t1 5.8005
R2699 a_11980_2192.n3 a_11980_2192.t3 5.8005
R2700 a_11980_2192.n3 a_11980_2192.t2 5.8005
R2701 a_11980_2192.n0 a_11980_2192.t7 5.8005
R2702 a_11980_2192.n0 a_11980_2192.t6 5.8005
R2703 a_11980_2192.t10 a_11980_2192.n10 5.8005
R2704 a_11980_2192.n10 a_11980_2192.t8 5.8005
R2705 a_11980_2192.n8 a_11980_2192.n6 1.94072
R2706 a_11980_2192.n9 a_11980_2192.n8 1.47876
R2707 a_11980_2192.n6 a_11980_2192.n5 0.478761
R2708 a_11980_2192.n5 a_11980_2192.n4 0.478761
R2709 saff_delay_unit_4/delay_unit_2_0.in_2.n8 saff_delay_unit_4/delay_unit_2_0.in_2.t14 784.053
R2710 saff_delay_unit_4/delay_unit_2_0.in_2.n8 saff_delay_unit_4/delay_unit_2_0.in_2.t10 784.053
R2711 saff_delay_unit_4/delay_unit_2_0.in_2.n9 saff_delay_unit_4/delay_unit_2_0.in_2.t12 784.053
R2712 saff_delay_unit_4/delay_unit_2_0.in_2.n9 saff_delay_unit_4/delay_unit_2_0.in_2.t16 784.053
R2713 saff_delay_unit_4/delay_unit_2_0.in_2.n3 saff_delay_unit_4/delay_unit_2_0.in_2.t18 523.774
R2714 saff_delay_unit_4/delay_unit_2_0.in_2.n4 saff_delay_unit_4/delay_unit_2_0.in_2.t9 523.774
R2715 saff_delay_unit_4/delay_unit_2_0.in_2.n0 saff_delay_unit_4/delay_unit_2_0.in_2.t17 523.774
R2716 saff_delay_unit_4/delay_unit_2_0.in_2.n1 saff_delay_unit_4/delay_unit_2_0.in_2.t11 523.774
R2717 saff_delay_unit_4/delay_unit_2_0.in_2.n3 saff_delay_unit_4/delay_unit_2_0.in_2.t8 202.44
R2718 saff_delay_unit_4/delay_unit_2_0.in_2.n4 saff_delay_unit_4/delay_unit_2_0.in_2.t13 202.44
R2719 saff_delay_unit_4/delay_unit_2_0.in_2.n0 saff_delay_unit_4/delay_unit_2_0.in_2.t19 202.44
R2720 saff_delay_unit_4/delay_unit_2_0.in_2.n1 saff_delay_unit_4/delay_unit_2_0.in_2.t15 202.44
R2721 saff_delay_unit_4/delay_unit_2_0.in_2.n10 saff_delay_unit_4/delay_unit_2_0.in_2.n8 168.659
R2722 saff_delay_unit_4/delay_unit_2_0.in_2.n10 saff_delay_unit_4/delay_unit_2_0.in_2.n9 167.992
R2723 saff_delay_unit_4/delay_unit_2_0.in_2.n6 saff_delay_unit_4/delay_unit_2_0.in_2.n2 166.144
R2724 saff_delay_unit_4/delay_unit_2_0.in_2.n6 saff_delay_unit_4/delay_unit_2_0.in_2.n5 165.8
R2725 saff_delay_unit_4/delay_unit_2_0.in_2.n7 saff_delay_unit_4/delay_unit_2_0.in_2.t7 85.2499
R2726 saff_delay_unit_4/delay_unit_2_0.in_2.n14 saff_delay_unit_4/delay_unit_2_0.in_2.t0 85.2499
R2727 saff_delay_unit_4/delay_unit_2_0.in_2.n14 saff_delay_unit_4/delay_unit_2_0.in_2.t4 83.7172
R2728 saff_delay_unit_4/delay_unit_2_0.in_2.n7 saff_delay_unit_4/delay_unit_2_0.in_2.t6 83.7172
R2729 saff_delay_unit_4/delay_unit_2_0.in_2.n13 saff_delay_unit_4/delay_unit_2_0.in_2.n11 75.7282
R2730 saff_delay_unit_4/delay_unit_2_0.in_2.n13 saff_delay_unit_4/delay_unit_2_0.in_2.n12 66.3172
R2731 saff_delay_unit_4/delay_unit_2_0.in_2.n5 saff_delay_unit_4/delay_unit_2_0.in_2.n3 27.8082
R2732 saff_delay_unit_4/delay_unit_2_0.in_2.n2 saff_delay_unit_4/delay_unit_2_0.in_2.n0 27.8082
R2733 saff_delay_unit_4/delay_unit_2_0.in_2.n5 saff_delay_unit_4/delay_unit_2_0.in_2.n4 26.5723
R2734 saff_delay_unit_4/delay_unit_2_0.in_2.n2 saff_delay_unit_4/delay_unit_2_0.in_2.n1 26.5723
R2735 saff_delay_unit_4/delay_unit_2_0.in_2.n12 saff_delay_unit_4/delay_unit_2_0.in_2.t1 17.4005
R2736 saff_delay_unit_4/delay_unit_2_0.in_2.n12 saff_delay_unit_4/delay_unit_2_0.in_2.t2 17.4005
R2737 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n10 17.1141
R2738 saff_delay_unit_4/delay_unit_2_0.in_2.n11 saff_delay_unit_4/delay_unit_2_0.in_2.t3 9.52217
R2739 saff_delay_unit_4/delay_unit_2_0.in_2.n11 saff_delay_unit_4/delay_unit_2_0.in_2.t5 9.52217
R2740 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n7 6.45821
R2741 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n13 5.30824
R2742 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n14 4.94887
R2743 saff_delay_unit_4/delay_unit_2_0.in_2.n15 saff_delay_unit_4/delay_unit_2_0.in_2 1.70362
R2744 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n6 1.06691
R2745 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2.n15 0.602062
R2746 saff_delay_unit_4/delay_unit_2_0.in_2.n15 saff_delay_unit_4/delay_unit_2_0.in_2 0.453625
R2747 saff_delay_unit_5/delay_unit_2_0.in_1.n13 saff_delay_unit_5/delay_unit_2_0.in_1.t18 572.12
R2748 saff_delay_unit_5/delay_unit_2_0.in_1.n13 saff_delay_unit_5/delay_unit_2_0.in_1.t12 572.12
R2749 saff_delay_unit_5/delay_unit_2_0.in_1.n12 saff_delay_unit_5/delay_unit_2_0.in_1.t10 572.12
R2750 saff_delay_unit_5/delay_unit_2_0.in_1.n12 saff_delay_unit_5/delay_unit_2_0.in_1.t14 572.12
R2751 saff_delay_unit_5/delay_unit_2_0.in_1.n3 saff_delay_unit_5/delay_unit_2_0.in_1.t17 523.774
R2752 saff_delay_unit_5/delay_unit_2_0.in_1.n4 saff_delay_unit_5/delay_unit_2_0.in_1.t11 523.774
R2753 saff_delay_unit_5/delay_unit_2_0.in_1.n0 saff_delay_unit_5/delay_unit_2_0.in_1.t19 523.774
R2754 saff_delay_unit_5/delay_unit_2_0.in_1.n1 saff_delay_unit_5/delay_unit_2_0.in_1.t13 523.774
R2755 saff_delay_unit_5/delay_unit_2_0.in_1.n3 saff_delay_unit_5/delay_unit_2_0.in_1.t8 202.44
R2756 saff_delay_unit_5/delay_unit_2_0.in_1.n4 saff_delay_unit_5/delay_unit_2_0.in_1.t15 202.44
R2757 saff_delay_unit_5/delay_unit_2_0.in_1.n0 saff_delay_unit_5/delay_unit_2_0.in_1.t9 202.44
R2758 saff_delay_unit_5/delay_unit_2_0.in_1.n1 saff_delay_unit_5/delay_unit_2_0.in_1.t16 202.44
R2759 saff_delay_unit_5/delay_unit_2_0.in_1.n14 saff_delay_unit_5/delay_unit_2_0.in_1.n12 166.468
R2760 saff_delay_unit_5/delay_unit_2_0.in_1.n6 saff_delay_unit_5/delay_unit_2_0.in_1.n2 166.149
R2761 saff_delay_unit_5/delay_unit_2_0.in_1.n14 saff_delay_unit_5/delay_unit_2_0.in_1.n13 165.8
R2762 saff_delay_unit_5/delay_unit_2_0.in_1.n6 saff_delay_unit_5/delay_unit_2_0.in_1.n5 165.8
R2763 saff_delay_unit_5/delay_unit_2_0.in_1.n7 saff_delay_unit_5/delay_unit_2_0.in_1.t0 85.1574
R2764 saff_delay_unit_5/delay_unit_2_0.in_1.n16 saff_delay_unit_5/delay_unit_2_0.in_1.t5 83.8097
R2765 saff_delay_unit_5/delay_unit_2_0.in_1.n7 saff_delay_unit_5/delay_unit_2_0.in_1.t7 83.8097
R2766 saff_delay_unit_5/delay_unit_2_0.in_1.n15 saff_delay_unit_5/delay_unit_2_0.in_1.t1 83.7172
R2767 saff_delay_unit_5/delay_unit_2_0.in_1.n11 saff_delay_unit_5/delay_unit_2_0.in_1.n10 74.288
R2768 saff_delay_unit_5/delay_unit_2_0.in_1.n11 saff_delay_unit_5/delay_unit_2_0.in_1.n9 67.7574
R2769 saff_delay_unit_5/delay_unit_2_0.in_1.n5 saff_delay_unit_5/delay_unit_2_0.in_1.n3 27.8082
R2770 saff_delay_unit_5/delay_unit_2_0.in_1.n2 saff_delay_unit_5/delay_unit_2_0.in_1.n1 27.8082
R2771 saff_delay_unit_5/delay_unit_2_0.in_1.n5 saff_delay_unit_5/delay_unit_2_0.in_1.n4 26.5723
R2772 saff_delay_unit_5/delay_unit_2_0.in_1.n2 saff_delay_unit_5/delay_unit_2_0.in_1.n0 26.5723
R2773 saff_delay_unit_5/delay_unit_2_0.in_1.n9 saff_delay_unit_5/delay_unit_2_0.in_1.t2 17.4005
R2774 saff_delay_unit_5/delay_unit_2_0.in_1.n9 saff_delay_unit_5/delay_unit_2_0.in_1.t3 17.4005
R2775 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_1.n14 16.0275
R2776 saff_delay_unit_5/delay_unit_2_0.in_1.n8 saff_delay_unit_5/delay_unit_2_0.in_1.n6 11.8364
R2777 saff_delay_unit_5/delay_unit_2_0.in_1.n10 saff_delay_unit_5/delay_unit_2_0.in_1.t6 9.52217
R2778 saff_delay_unit_5/delay_unit_2_0.in_1.n10 saff_delay_unit_5/delay_unit_2_0.in_1.t4 9.52217
R2779 saff_delay_unit_5/delay_unit_2_0.in_1.n15 saff_delay_unit_5/delay_unit_2_0.in_1 6.02878
R2780 saff_delay_unit_5/delay_unit_2_0.in_1.n17 saff_delay_unit_5/delay_unit_2_0.in_1.n11 5.83219
R2781 saff_delay_unit_5/delay_unit_2_0.in_1.n8 saff_delay_unit_5/delay_unit_2_0.in_1.n7 5.74235
R2782 saff_delay_unit_5/delay_unit_2_0.in_1.n17 saff_delay_unit_5/delay_unit_2_0.in_1.n16 5.49235
R2783 saff_delay_unit_5/delay_unit_2_0.in_1.n16 saff_delay_unit_5/delay_unit_2_0.in_1.n15 1.44072
R2784 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_1.n17 1.32081
R2785 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_1.n8 0.285656
R2786 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 879.481
R2787 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 742.783
R2788 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 665.16
R2789 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 623.388
R2790 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 523.774
R2791 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 431.807
R2792 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 427.875
R2793 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 357.26
R2794 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 208.537
R2795 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 168.077
R2796 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R2797 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R2798 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R2799 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 11.1806
R2800 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R2801 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R2802 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R2803 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R2804 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R2805 saff_delay_unit_2/delay_unit_2_0.in_1.n12 saff_delay_unit_2/delay_unit_2_0.in_1.t16 572.12
R2806 saff_delay_unit_2/delay_unit_2_0.in_1.n12 saff_delay_unit_2/delay_unit_2_0.in_1.t9 572.12
R2807 saff_delay_unit_2/delay_unit_2_0.in_1.n11 saff_delay_unit_2/delay_unit_2_0.in_1.t13 572.12
R2808 saff_delay_unit_2/delay_unit_2_0.in_1.n11 saff_delay_unit_2/delay_unit_2_0.in_1.t18 572.12
R2809 saff_delay_unit_2/delay_unit_2_0.in_1.n3 saff_delay_unit_2/delay_unit_2_0.in_1.t19 523.774
R2810 saff_delay_unit_2/delay_unit_2_0.in_1.n4 saff_delay_unit_2/delay_unit_2_0.in_1.t12 523.774
R2811 saff_delay_unit_2/delay_unit_2_0.in_1.n0 saff_delay_unit_2/delay_unit_2_0.in_1.t8 523.774
R2812 saff_delay_unit_2/delay_unit_2_0.in_1.n1 saff_delay_unit_2/delay_unit_2_0.in_1.t14 523.774
R2813 saff_delay_unit_2/delay_unit_2_0.in_1.n3 saff_delay_unit_2/delay_unit_2_0.in_1.t10 202.44
R2814 saff_delay_unit_2/delay_unit_2_0.in_1.n4 saff_delay_unit_2/delay_unit_2_0.in_1.t15 202.44
R2815 saff_delay_unit_2/delay_unit_2_0.in_1.n0 saff_delay_unit_2/delay_unit_2_0.in_1.t11 202.44
R2816 saff_delay_unit_2/delay_unit_2_0.in_1.n1 saff_delay_unit_2/delay_unit_2_0.in_1.t17 202.44
R2817 saff_delay_unit_2/delay_unit_2_0.in_1.n13 saff_delay_unit_2/delay_unit_2_0.in_1.n11 166.468
R2818 saff_delay_unit_2/delay_unit_2_0.in_1.n6 saff_delay_unit_2/delay_unit_2_0.in_1.n2 166.149
R2819 saff_delay_unit_2/delay_unit_2_0.in_1.n6 saff_delay_unit_2/delay_unit_2_0.in_1.n5 165.8
R2820 saff_delay_unit_2/delay_unit_2_0.in_1.n13 saff_delay_unit_2/delay_unit_2_0.in_1.n12 165.8
R2821 saff_delay_unit_2/delay_unit_2_0.in_1.n7 saff_delay_unit_2/delay_unit_2_0.in_1.t0 85.1574
R2822 saff_delay_unit_2/delay_unit_2_0.in_1.n15 saff_delay_unit_2/delay_unit_2_0.in_1.t4 83.8097
R2823 saff_delay_unit_2/delay_unit_2_0.in_1.n7 saff_delay_unit_2/delay_unit_2_0.in_1.t1 83.8097
R2824 saff_delay_unit_2/delay_unit_2_0.in_1.n14 saff_delay_unit_2/delay_unit_2_0.in_1.t5 83.7172
R2825 saff_delay_unit_2/delay_unit_2_0.in_1.n10 saff_delay_unit_2/delay_unit_2_0.in_1.n9 74.288
R2826 saff_delay_unit_2/delay_unit_2_0.in_1.n10 saff_delay_unit_2/delay_unit_2_0.in_1.n8 67.7574
R2827 saff_delay_unit_2/delay_unit_2_0.in_1.n5 saff_delay_unit_2/delay_unit_2_0.in_1.n3 27.8082
R2828 saff_delay_unit_2/delay_unit_2_0.in_1.n2 saff_delay_unit_2/delay_unit_2_0.in_1.n1 27.8082
R2829 saff_delay_unit_2/delay_unit_2_0.in_1.n5 saff_delay_unit_2/delay_unit_2_0.in_1.n4 26.5723
R2830 saff_delay_unit_2/delay_unit_2_0.in_1.n2 saff_delay_unit_2/delay_unit_2_0.in_1.n0 26.5723
R2831 saff_delay_unit_2/delay_unit_2_0.in_1.n8 saff_delay_unit_2/delay_unit_2_0.in_1.t6 17.4005
R2832 saff_delay_unit_2/delay_unit_2_0.in_1.n8 saff_delay_unit_2/delay_unit_2_0.in_1.t2 17.4005
R2833 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/delay_unit_2_0.in_1.n13 16.0275
R2834 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/delay_unit_2_0.in_1.n6 11.8364
R2835 saff_delay_unit_2/delay_unit_2_0.in_1.n9 saff_delay_unit_2/delay_unit_2_0.in_1.t3 9.52217
R2836 saff_delay_unit_2/delay_unit_2_0.in_1.n9 saff_delay_unit_2/delay_unit_2_0.in_1.t7 9.52217
R2837 saff_delay_unit_2/delay_unit_2_0.in_1.n14 saff_delay_unit_2/delay_unit_2_0.in_1 6.02878
R2838 saff_delay_unit_2/delay_unit_2_0.in_1.n16 saff_delay_unit_2/delay_unit_2_0.in_1.n10 5.83219
R2839 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/delay_unit_2_0.in_1.n7 5.74235
R2840 saff_delay_unit_2/delay_unit_2_0.in_1.n16 saff_delay_unit_2/delay_unit_2_0.in_1.n15 5.49235
R2841 saff_delay_unit_2/delay_unit_2_0.in_1.n15 saff_delay_unit_2/delay_unit_2_0.in_1.n14 1.44072
R2842 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/delay_unit_2_0.in_1.n16 1.32081
R2843 saff_delay_unit_3/delay_unit_2_0.in_2.n8 saff_delay_unit_3/delay_unit_2_0.in_2.t11 784.053
R2844 saff_delay_unit_3/delay_unit_2_0.in_2.n8 saff_delay_unit_3/delay_unit_2_0.in_2.t16 784.053
R2845 saff_delay_unit_3/delay_unit_2_0.in_2.n9 saff_delay_unit_3/delay_unit_2_0.in_2.t12 784.053
R2846 saff_delay_unit_3/delay_unit_2_0.in_2.n9 saff_delay_unit_3/delay_unit_2_0.in_2.t8 784.053
R2847 saff_delay_unit_3/delay_unit_2_0.in_2.n3 saff_delay_unit_3/delay_unit_2_0.in_2.t14 523.774
R2848 saff_delay_unit_3/delay_unit_2_0.in_2.n4 saff_delay_unit_3/delay_unit_2_0.in_2.t19 523.774
R2849 saff_delay_unit_3/delay_unit_2_0.in_2.n0 saff_delay_unit_3/delay_unit_2_0.in_2.t13 523.774
R2850 saff_delay_unit_3/delay_unit_2_0.in_2.n1 saff_delay_unit_3/delay_unit_2_0.in_2.t18 523.774
R2851 saff_delay_unit_3/delay_unit_2_0.in_2.n3 saff_delay_unit_3/delay_unit_2_0.in_2.t17 202.44
R2852 saff_delay_unit_3/delay_unit_2_0.in_2.n4 saff_delay_unit_3/delay_unit_2_0.in_2.t10 202.44
R2853 saff_delay_unit_3/delay_unit_2_0.in_2.n0 saff_delay_unit_3/delay_unit_2_0.in_2.t15 202.44
R2854 saff_delay_unit_3/delay_unit_2_0.in_2.n1 saff_delay_unit_3/delay_unit_2_0.in_2.t9 202.44
R2855 saff_delay_unit_3/delay_unit_2_0.in_2.n10 saff_delay_unit_3/delay_unit_2_0.in_2.n8 168.659
R2856 saff_delay_unit_3/delay_unit_2_0.in_2.n10 saff_delay_unit_3/delay_unit_2_0.in_2.n9 167.992
R2857 saff_delay_unit_3/delay_unit_2_0.in_2.n6 saff_delay_unit_3/delay_unit_2_0.in_2.n2 166.144
R2858 saff_delay_unit_3/delay_unit_2_0.in_2.n6 saff_delay_unit_3/delay_unit_2_0.in_2.n5 165.8
R2859 saff_delay_unit_3/delay_unit_2_0.in_2.n7 saff_delay_unit_3/delay_unit_2_0.in_2.t6 85.2499
R2860 saff_delay_unit_3/delay_unit_2_0.in_2.n14 saff_delay_unit_3/delay_unit_2_0.in_2.t5 85.2499
R2861 saff_delay_unit_3/delay_unit_2_0.in_2.n14 saff_delay_unit_3/delay_unit_2_0.in_2.t1 83.7172
R2862 saff_delay_unit_3/delay_unit_2_0.in_2.n7 saff_delay_unit_3/delay_unit_2_0.in_2.t7 83.7172
R2863 saff_delay_unit_3/delay_unit_2_0.in_2.n13 saff_delay_unit_3/delay_unit_2_0.in_2.n11 75.7282
R2864 saff_delay_unit_3/delay_unit_2_0.in_2.n13 saff_delay_unit_3/delay_unit_2_0.in_2.n12 66.3172
R2865 saff_delay_unit_3/delay_unit_2_0.in_2.n5 saff_delay_unit_3/delay_unit_2_0.in_2.n3 27.8082
R2866 saff_delay_unit_3/delay_unit_2_0.in_2.n2 saff_delay_unit_3/delay_unit_2_0.in_2.n0 27.8082
R2867 saff_delay_unit_3/delay_unit_2_0.in_2.n5 saff_delay_unit_3/delay_unit_2_0.in_2.n4 26.5723
R2868 saff_delay_unit_3/delay_unit_2_0.in_2.n2 saff_delay_unit_3/delay_unit_2_0.in_2.n1 26.5723
R2869 saff_delay_unit_3/delay_unit_2_0.in_2.n12 saff_delay_unit_3/delay_unit_2_0.in_2.t0 17.4005
R2870 saff_delay_unit_3/delay_unit_2_0.in_2.n12 saff_delay_unit_3/delay_unit_2_0.in_2.t2 17.4005
R2871 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2.n10 17.1141
R2872 saff_delay_unit_3/delay_unit_2_0.in_2.n11 saff_delay_unit_3/delay_unit_2_0.in_2.t4 9.52217
R2873 saff_delay_unit_3/delay_unit_2_0.in_2.n11 saff_delay_unit_3/delay_unit_2_0.in_2.t3 9.52217
R2874 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2.n7 6.45821
R2875 saff_delay_unit_3/delay_unit_2_0.in_2.n15 saff_delay_unit_3/delay_unit_2_0.in_2.n13 5.30824
R2876 saff_delay_unit_3/delay_unit_2_0.in_2.n15 saff_delay_unit_3/delay_unit_2_0.in_2.n14 4.94887
R2877 saff_delay_unit_3/delay_unit_2_0.in_2.n16 saff_delay_unit_3/delay_unit_2_0.in_2 1.54347
R2878 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2.n6 1.06691
R2879 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2.n16 0.602062
R2880 saff_delay_unit_3/delay_unit_2_0.in_2.n16 saff_delay_unit_3/delay_unit_2_0.in_2 0.453625
R2881 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2.n15 0.160656
R2882 start_pos.n3 start_pos.t5 523.774
R2883 start_pos.n4 start_pos.t7 523.774
R2884 start_pos.n0 start_pos.t4 523.774
R2885 start_pos.n1 start_pos.t9 523.774
R2886 start_pos.n3 start_pos.t8 202.44
R2887 start_pos.n4 start_pos.t2 202.44
R2888 start_pos.n0 start_pos.t6 202.44
R2889 start_pos.n1 start_pos.t3 202.44
R2890 start_pos.n6 start_pos.n2 166.149
R2891 start_pos.n6 start_pos.n5 165.8
R2892 start_pos.n7 start_pos.t1 85.1574
R2893 start_pos.n7 start_pos.t0 83.8097
R2894 start_pos.n5 start_pos.n3 27.8082
R2895 start_pos.n2 start_pos.n1 27.8082
R2896 start_pos.n5 start_pos.n4 26.5723
R2897 start_pos.n2 start_pos.n0 26.5723
R2898 start_pos.n8 start_pos.n6 11.8364
R2899 start_pos.n8 start_pos.n7 5.74235
R2900 start_pos start_pos.n8 0.285656
R2901 start_neg.n4 start_neg.t5 523.774
R2902 start_neg.n5 start_neg.t9 523.774
R2903 start_neg.n1 start_neg.t6 523.774
R2904 start_neg.n2 start_neg.t2 523.774
R2905 start_neg.n4 start_neg.t7 202.44
R2906 start_neg.n5 start_neg.t3 202.44
R2907 start_neg.n1 start_neg.t8 202.44
R2908 start_neg.n2 start_neg.t4 202.44
R2909 start_neg.n7 start_neg.n3 166.144
R2910 start_neg.n7 start_neg.n6 165.8
R2911 start_neg.n0 start_neg.t1 85.2499
R2912 start_neg.n0 start_neg.t0 83.7172
R2913 start_neg.n6 start_neg.n4 27.8082
R2914 start_neg.n3 start_neg.n1 27.8082
R2915 start_neg.n6 start_neg.n5 26.5723
R2916 start_neg.n3 start_neg.n2 26.5723
R2917 start_neg.n8 start_neg.n0 6.45821
R2918 start_neg start_neg.n7 0.879406
R2919 start_neg.n8 start_neg 0.188
R2920 start_neg start_neg.n8 0.063
R2921 saff_delay_unit_1/delay_unit_2_0.in_2.n8 saff_delay_unit_1/delay_unit_2_0.in_2.t10 784.053
R2922 saff_delay_unit_1/delay_unit_2_0.in_2.n8 saff_delay_unit_1/delay_unit_2_0.in_2.t13 784.053
R2923 saff_delay_unit_1/delay_unit_2_0.in_2.n9 saff_delay_unit_1/delay_unit_2_0.in_2.t9 784.053
R2924 saff_delay_unit_1/delay_unit_2_0.in_2.n9 saff_delay_unit_1/delay_unit_2_0.in_2.t15 784.053
R2925 saff_delay_unit_1/delay_unit_2_0.in_2.n3 saff_delay_unit_1/delay_unit_2_0.in_2.t14 523.774
R2926 saff_delay_unit_1/delay_unit_2_0.in_2.n4 saff_delay_unit_1/delay_unit_2_0.in_2.t18 523.774
R2927 saff_delay_unit_1/delay_unit_2_0.in_2.n0 saff_delay_unit_1/delay_unit_2_0.in_2.t17 523.774
R2928 saff_delay_unit_1/delay_unit_2_0.in_2.n1 saff_delay_unit_1/delay_unit_2_0.in_2.t19 523.774
R2929 saff_delay_unit_1/delay_unit_2_0.in_2.n3 saff_delay_unit_1/delay_unit_2_0.in_2.t16 202.44
R2930 saff_delay_unit_1/delay_unit_2_0.in_2.n4 saff_delay_unit_1/delay_unit_2_0.in_2.t11 202.44
R2931 saff_delay_unit_1/delay_unit_2_0.in_2.n0 saff_delay_unit_1/delay_unit_2_0.in_2.t8 202.44
R2932 saff_delay_unit_1/delay_unit_2_0.in_2.n1 saff_delay_unit_1/delay_unit_2_0.in_2.t12 202.44
R2933 saff_delay_unit_1/delay_unit_2_0.in_2.n10 saff_delay_unit_1/delay_unit_2_0.in_2.n8 168.659
R2934 saff_delay_unit_1/delay_unit_2_0.in_2.n10 saff_delay_unit_1/delay_unit_2_0.in_2.n9 167.992
R2935 saff_delay_unit_1/delay_unit_2_0.in_2.n6 saff_delay_unit_1/delay_unit_2_0.in_2.n2 166.144
R2936 saff_delay_unit_1/delay_unit_2_0.in_2.n6 saff_delay_unit_1/delay_unit_2_0.in_2.n5 165.8
R2937 saff_delay_unit_1/delay_unit_2_0.in_2.n7 saff_delay_unit_1/delay_unit_2_0.in_2.t1 85.2499
R2938 saff_delay_unit_1/delay_unit_2_0.in_2.n14 saff_delay_unit_1/delay_unit_2_0.in_2.t7 85.2499
R2939 saff_delay_unit_1/delay_unit_2_0.in_2.n14 saff_delay_unit_1/delay_unit_2_0.in_2.t3 83.7172
R2940 saff_delay_unit_1/delay_unit_2_0.in_2.n7 saff_delay_unit_1/delay_unit_2_0.in_2.t0 83.7172
R2941 saff_delay_unit_1/delay_unit_2_0.in_2.n13 saff_delay_unit_1/delay_unit_2_0.in_2.n11 75.7282
R2942 saff_delay_unit_1/delay_unit_2_0.in_2.n13 saff_delay_unit_1/delay_unit_2_0.in_2.n12 66.3172
R2943 saff_delay_unit_1/delay_unit_2_0.in_2.n5 saff_delay_unit_1/delay_unit_2_0.in_2.n3 27.8082
R2944 saff_delay_unit_1/delay_unit_2_0.in_2.n2 saff_delay_unit_1/delay_unit_2_0.in_2.n0 27.8082
R2945 saff_delay_unit_1/delay_unit_2_0.in_2.n5 saff_delay_unit_1/delay_unit_2_0.in_2.n4 26.5723
R2946 saff_delay_unit_1/delay_unit_2_0.in_2.n2 saff_delay_unit_1/delay_unit_2_0.in_2.n1 26.5723
R2947 saff_delay_unit_1/delay_unit_2_0.in_2.n12 saff_delay_unit_1/delay_unit_2_0.in_2.t4 17.4005
R2948 saff_delay_unit_1/delay_unit_2_0.in_2.n12 saff_delay_unit_1/delay_unit_2_0.in_2.t2 17.4005
R2949 saff_delay_unit_1/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2.n10 17.1141
R2950 saff_delay_unit_1/delay_unit_2_0.in_2.n11 saff_delay_unit_1/delay_unit_2_0.in_2.t5 9.52217
R2951 saff_delay_unit_1/delay_unit_2_0.in_2.n11 saff_delay_unit_1/delay_unit_2_0.in_2.t6 9.52217
R2952 saff_delay_unit_1/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2.n7 6.45821
R2953 saff_delay_unit_1/delay_unit_2_0.in_2.n15 saff_delay_unit_1/delay_unit_2_0.in_2.n13 5.30824
R2954 saff_delay_unit_1/delay_unit_2_0.in_2.n15 saff_delay_unit_1/delay_unit_2_0.in_2.n14 4.94887
R2955 saff_delay_unit_1/delay_unit_2_0.in_2.n16 saff_delay_unit_1/delay_unit_2_0.in_2 1.54347
R2956 saff_delay_unit_1/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2.n6 1.06691
R2957 saff_delay_unit_1/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2.n16 0.602062
R2958 saff_delay_unit_1/delay_unit_2_0.in_2.n16 saff_delay_unit_1/delay_unit_2_0.in_2 0.453625
R2959 saff_delay_unit_1/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2.n15 0.160656
R2960 a_834_2192.n2 a_834_2192.n1 34.9195
R2961 a_834_2192.n3 a_834_2192.n2 25.5407
R2962 a_834_2192.n2 a_834_2192.n0 25.2907
R2963 a_834_2192.n1 a_834_2192.t4 5.8005
R2964 a_834_2192.n1 a_834_2192.t3 5.8005
R2965 a_834_2192.n0 a_834_2192.t5 5.8005
R2966 a_834_2192.n0 a_834_2192.t2 5.8005
R2967 a_834_2192.n3 a_834_2192.t1 5.8005
R2968 a_834_2192.t0 a_834_2192.n3 5.8005
R2969 a_570_2192.n4 a_570_2192.t2 32.0282
R2970 a_570_2192.n9 a_570_2192.n0 25.7663
R2971 a_570_2192.n6 a_570_2192.n1 25.75
R2972 a_570_2192.n5 a_570_2192.n2 25.75
R2973 a_570_2192.n4 a_570_2192.n3 25.75
R2974 a_570_2192.n10 a_570_2192.n9 25.288
R2975 a_570_2192.n8 a_570_2192.n7 24.288
R2976 a_570_2192.n7 a_570_2192.t5 5.8005
R2977 a_570_2192.n7 a_570_2192.t12 5.8005
R2978 a_570_2192.n1 a_570_2192.t9 5.8005
R2979 a_570_2192.n1 a_570_2192.t0 5.8005
R2980 a_570_2192.n2 a_570_2192.t3 5.8005
R2981 a_570_2192.n2 a_570_2192.t11 5.8005
R2982 a_570_2192.n3 a_570_2192.t10 5.8005
R2983 a_570_2192.n3 a_570_2192.t1 5.8005
R2984 a_570_2192.n0 a_570_2192.t4 5.8005
R2985 a_570_2192.n0 a_570_2192.t7 5.8005
R2986 a_570_2192.n10 a_570_2192.t6 5.8005
R2987 a_570_2192.t8 a_570_2192.n10 5.8005
R2988 a_570_2192.n8 a_570_2192.n6 1.94072
R2989 a_570_2192.n9 a_570_2192.n8 1.47876
R2990 a_570_2192.n6 a_570_2192.n5 0.478761
R2991 a_570_2192.n5 a_570_2192.n4 0.478761
R2992 saff_delay_unit_7/saff_2_0.d.n12 saff_delay_unit_7/saff_2_0.d.t8 572.12
R2993 saff_delay_unit_7/saff_2_0.d.n12 saff_delay_unit_7/saff_2_0.d.t10 572.12
R2994 saff_delay_unit_7/saff_2_0.d.n11 saff_delay_unit_7/saff_2_0.d.t14 572.12
R2995 saff_delay_unit_7/saff_2_0.d.n11 saff_delay_unit_7/saff_2_0.d.t15 572.12
R2996 saff_delay_unit_7/saff_2_0.d.n3 saff_delay_unit_7/saff_2_0.d.t19 523.774
R2997 saff_delay_unit_7/saff_2_0.d.n4 saff_delay_unit_7/saff_2_0.d.t13 523.774
R2998 saff_delay_unit_7/saff_2_0.d.n0 saff_delay_unit_7/saff_2_0.d.t9 523.774
R2999 saff_delay_unit_7/saff_2_0.d.n1 saff_delay_unit_7/saff_2_0.d.t16 523.774
R3000 saff_delay_unit_7/saff_2_0.d.n3 saff_delay_unit_7/saff_2_0.d.t11 202.44
R3001 saff_delay_unit_7/saff_2_0.d.n4 saff_delay_unit_7/saff_2_0.d.t17 202.44
R3002 saff_delay_unit_7/saff_2_0.d.n0 saff_delay_unit_7/saff_2_0.d.t12 202.44
R3003 saff_delay_unit_7/saff_2_0.d.n1 saff_delay_unit_7/saff_2_0.d.t18 202.44
R3004 saff_delay_unit_7/saff_2_0.d.n13 saff_delay_unit_7/saff_2_0.d.n11 166.468
R3005 saff_delay_unit_7/saff_2_0.d.n6 saff_delay_unit_7/saff_2_0.d.n2 166.149
R3006 saff_delay_unit_7/saff_2_0.d.n13 saff_delay_unit_7/saff_2_0.d.n12 165.8
R3007 saff_delay_unit_7/saff_2_0.d.n6 saff_delay_unit_7/saff_2_0.d.n5 165.8
R3008 saff_delay_unit_7/saff_2_0.d.n7 saff_delay_unit_7/saff_2_0.d.t0 85.1574
R3009 saff_delay_unit_7/saff_2_0.d.n15 saff_delay_unit_7/saff_2_0.d.t6 83.8097
R3010 saff_delay_unit_7/saff_2_0.d.n7 saff_delay_unit_7/saff_2_0.d.t2 83.8097
R3011 saff_delay_unit_7/saff_2_0.d.n14 saff_delay_unit_7/saff_2_0.d.t3 83.7172
R3012 saff_delay_unit_7/saff_2_0.d.n10 saff_delay_unit_7/saff_2_0.d.n9 74.288
R3013 saff_delay_unit_7/saff_2_0.d.n10 saff_delay_unit_7/saff_2_0.d.n8 67.7574
R3014 saff_delay_unit_7/saff_2_0.d.n5 saff_delay_unit_7/saff_2_0.d.n3 27.8082
R3015 saff_delay_unit_7/saff_2_0.d.n2 saff_delay_unit_7/saff_2_0.d.n1 27.8082
R3016 saff_delay_unit_7/saff_2_0.d.n5 saff_delay_unit_7/saff_2_0.d.n4 26.5723
R3017 saff_delay_unit_7/saff_2_0.d.n2 saff_delay_unit_7/saff_2_0.d.n0 26.5723
R3018 saff_delay_unit_7/saff_2_0.d.n8 saff_delay_unit_7/saff_2_0.d.t7 17.4005
R3019 saff_delay_unit_7/saff_2_0.d.n8 saff_delay_unit_7/saff_2_0.d.t4 17.4005
R3020 saff_delay_unit_7/saff_2_0.sense_amplifier_0.d saff_delay_unit_7/saff_2_0.d.n13 16.0275
R3021 delay_unit_2_0.in_1 saff_delay_unit_7/saff_2_0.d.n6 11.8364
R3022 saff_delay_unit_7/saff_2_0.d.n9 saff_delay_unit_7/saff_2_0.d.t5 9.52217
R3023 saff_delay_unit_7/saff_2_0.d.n9 saff_delay_unit_7/saff_2_0.d.t1 9.52217
R3024 saff_delay_unit_7/saff_2_0.d.n14 saff_delay_unit_7/saff_2_0.sense_amplifier_0.d 6.02878
R3025 saff_delay_unit_7/saff_2_0.d.n16 saff_delay_unit_7/saff_2_0.d.n10 5.83219
R3026 delay_unit_2_0.in_1 saff_delay_unit_7/saff_2_0.d.n7 5.74235
R3027 saff_delay_unit_7/saff_2_0.d.n16 saff_delay_unit_7/saff_2_0.d.n15 5.49235
R3028 saff_delay_unit_7/delay_unit_2_0.out_1 delay_unit_2_0.in_1 2.48878
R3029 saff_delay_unit_7/saff_2_0.d.n15 saff_delay_unit_7/saff_2_0.d.n14 1.44072
R3030 saff_delay_unit_7/delay_unit_2_0.out_1 saff_delay_unit_7/saff_2_0.d.n16 1.32081
R3031 a_16544_2192.n4 a_16544_2192.t11 32.0282
R3032 a_16544_2192.n10 a_16544_2192.n9 25.7663
R3033 a_16544_2192.n6 a_16544_2192.n1 25.75
R3034 a_16544_2192.n5 a_16544_2192.n2 25.75
R3035 a_16544_2192.n4 a_16544_2192.n3 25.75
R3036 a_16544_2192.n9 a_16544_2192.n0 25.288
R3037 a_16544_2192.n8 a_16544_2192.n7 24.288
R3038 a_16544_2192.n7 a_16544_2192.t4 5.8005
R3039 a_16544_2192.n7 a_16544_2192.t2 5.8005
R3040 a_16544_2192.n1 a_16544_2192.t0 5.8005
R3041 a_16544_2192.n1 a_16544_2192.t10 5.8005
R3042 a_16544_2192.n2 a_16544_2192.t9 5.8005
R3043 a_16544_2192.n2 a_16544_2192.t3 5.8005
R3044 a_16544_2192.n3 a_16544_2192.t1 5.8005
R3045 a_16544_2192.n3 a_16544_2192.t12 5.8005
R3046 a_16544_2192.n0 a_16544_2192.t7 5.8005
R3047 a_16544_2192.n0 a_16544_2192.t6 5.8005
R3048 a_16544_2192.t8 a_16544_2192.n10 5.8005
R3049 a_16544_2192.n10 a_16544_2192.t5 5.8005
R3050 a_16544_2192.n8 a_16544_2192.n6 1.94072
R3051 a_16544_2192.n9 a_16544_2192.n8 1.47876
R3052 a_16544_2192.n6 a_16544_2192.n5 0.478761
R3053 a_16544_2192.n5 a_16544_2192.n4 0.478761
R3054 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 890.727
R3055 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 742.783
R3056 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 665.16
R3057 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 623.388
R3058 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 523.774
R3059 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 431.807
R3060 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 427.875
R3061 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 364.733
R3062 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 208.5
R3063 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 168.007
R3064 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R3065 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 31.2728
R3066 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 31.0337
R3067 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R3068 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R3069 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R3070 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 8.00471
R3071 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R3072 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3073 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R3074 term_3.n1 term_3.t5 734.539
R3075 term_3.n1 term_3.t4 233.26
R3076 term_3.n2 term_3.n1 162.399
R3077 term_3.n2 term_3.n0 75.5108
R3078 term_3.n4 term_3.n3 66.3172
R3079 term_3.n3 term_3.t2 17.4005
R3080 term_3.n3 term_3.t0 17.4005
R3081 term_3.n0 term_3.t1 9.52217
R3082 term_3.n0 term_3.t3 9.52217
R3083 term_3 term_3.n4 5.08746
R3084 term_3.n4 term_3.n2 0.3755
R3085 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 879.481
R3086 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 742.783
R3087 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 665.16
R3088 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 623.388
R3089 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 523.774
R3090 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 431.807
R3091 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 427.875
R3092 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 357.26
R3093 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 208.537
R3094 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 168.077
R3095 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R3096 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 31.2347
R3097 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R3098 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 11.1806
R3099 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R3100 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R3101 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R3102 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R3103 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R3104 saff_delay_unit_7/delay_unit_2_0.in_1.n1 saff_delay_unit_7/delay_unit_2_0.in_1.t13 572.12
R3105 saff_delay_unit_7/delay_unit_2_0.in_1.n1 saff_delay_unit_7/delay_unit_2_0.in_1.t8 572.12
R3106 saff_delay_unit_7/delay_unit_2_0.in_1.n0 saff_delay_unit_7/delay_unit_2_0.in_1.t17 572.12
R3107 saff_delay_unit_7/delay_unit_2_0.in_1.n0 saff_delay_unit_7/delay_unit_2_0.in_1.t12 572.12
R3108 saff_delay_unit_7/delay_unit_2_0.in_1.n6 saff_delay_unit_7/delay_unit_2_0.in_1.t14 523.774
R3109 saff_delay_unit_7/delay_unit_2_0.in_1.n7 saff_delay_unit_7/delay_unit_2_0.in_1.t16 523.774
R3110 saff_delay_unit_7/delay_unit_2_0.in_1.n3 saff_delay_unit_7/delay_unit_2_0.in_1.t18 523.774
R3111 saff_delay_unit_7/delay_unit_2_0.in_1.n4 saff_delay_unit_7/delay_unit_2_0.in_1.t19 523.774
R3112 saff_delay_unit_7/delay_unit_2_0.in_1.n6 saff_delay_unit_7/delay_unit_2_0.in_1.t15 202.44
R3113 saff_delay_unit_7/delay_unit_2_0.in_1.n7 saff_delay_unit_7/delay_unit_2_0.in_1.t9 202.44
R3114 saff_delay_unit_7/delay_unit_2_0.in_1.n3 saff_delay_unit_7/delay_unit_2_0.in_1.t10 202.44
R3115 saff_delay_unit_7/delay_unit_2_0.in_1.n4 saff_delay_unit_7/delay_unit_2_0.in_1.t11 202.44
R3116 saff_delay_unit_7/delay_unit_2_0.in_1.n2 saff_delay_unit_7/delay_unit_2_0.in_1.n0 166.468
R3117 saff_delay_unit_7/delay_unit_2_0.in_1.n9 saff_delay_unit_7/delay_unit_2_0.in_1.n5 166.149
R3118 saff_delay_unit_7/delay_unit_2_0.in_1.n9 saff_delay_unit_7/delay_unit_2_0.in_1.n8 165.8
R3119 saff_delay_unit_7/delay_unit_2_0.in_1.n2 saff_delay_unit_7/delay_unit_2_0.in_1.n1 165.8
R3120 saff_delay_unit_7/delay_unit_2_0.in_1.n10 saff_delay_unit_7/delay_unit_2_0.in_1.t1 85.1574
R3121 saff_delay_unit_7/delay_unit_2_0.in_1.n10 saff_delay_unit_7/delay_unit_2_0.in_1.t4 83.8097
R3122 saff_delay_unit_7/delay_unit_2_0.in_1.n15 saff_delay_unit_7/delay_unit_2_0.in_1.t2 83.8097
R3123 saff_delay_unit_7/delay_unit_2_0.in_1.n16 saff_delay_unit_7/delay_unit_2_0.in_1.t5 83.7172
R3124 saff_delay_unit_7/delay_unit_2_0.in_1.n13 saff_delay_unit_7/delay_unit_2_0.in_1.n12 74.288
R3125 saff_delay_unit_7/delay_unit_2_0.in_1.n13 saff_delay_unit_7/delay_unit_2_0.in_1.n11 67.7574
R3126 saff_delay_unit_7/delay_unit_2_0.in_1.n8 saff_delay_unit_7/delay_unit_2_0.in_1.n6 27.8082
R3127 saff_delay_unit_7/delay_unit_2_0.in_1.n5 saff_delay_unit_7/delay_unit_2_0.in_1.n4 27.8082
R3128 saff_delay_unit_7/delay_unit_2_0.in_1.n8 saff_delay_unit_7/delay_unit_2_0.in_1.n7 26.5723
R3129 saff_delay_unit_7/delay_unit_2_0.in_1.n5 saff_delay_unit_7/delay_unit_2_0.in_1.n3 26.5723
R3130 saff_delay_unit_7/delay_unit_2_0.in_1.n11 saff_delay_unit_7/delay_unit_2_0.in_1.t0 17.4005
R3131 saff_delay_unit_7/delay_unit_2_0.in_1.n11 saff_delay_unit_7/delay_unit_2_0.in_1.t7 17.4005
R3132 saff_delay_unit_7/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_1.n2 16.0275
R3133 saff_delay_unit_7/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_1.n9 11.8364
R3134 saff_delay_unit_7/delay_unit_2_0.in_1.n12 saff_delay_unit_7/delay_unit_2_0.in_1.t3 9.52217
R3135 saff_delay_unit_7/delay_unit_2_0.in_1.n12 saff_delay_unit_7/delay_unit_2_0.in_1.t6 9.52217
R3136 saff_delay_unit_7/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_1.n16 6.02878
R3137 saff_delay_unit_7/delay_unit_2_0.in_1.n14 saff_delay_unit_7/delay_unit_2_0.in_1.n13 5.83219
R3138 saff_delay_unit_7/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_1.n10 5.74235
R3139 saff_delay_unit_7/delay_unit_2_0.in_1.n15 saff_delay_unit_7/delay_unit_2_0.in_1.n14 5.49235
R3140 saff_delay_unit_7/delay_unit_2_0.in_1.n16 saff_delay_unit_7/delay_unit_2_0.in_1.n15 1.44072
R3141 saff_delay_unit_7/delay_unit_2_0.in_1.n14 saff_delay_unit_7/delay_unit_2_0.in_1 1.32081
R3142 a_14262_2192.n4 a_14262_2192.t3 32.0282
R3143 a_14262_2192.n10 a_14262_2192.n9 25.7663
R3144 a_14262_2192.n6 a_14262_2192.n1 25.75
R3145 a_14262_2192.n5 a_14262_2192.n2 25.75
R3146 a_14262_2192.n4 a_14262_2192.n3 25.75
R3147 a_14262_2192.n9 a_14262_2192.n0 25.288
R3148 a_14262_2192.n8 a_14262_2192.n7 24.288
R3149 a_14262_2192.n7 a_14262_2192.t10 5.8005
R3150 a_14262_2192.n7 a_14262_2192.t6 5.8005
R3151 a_14262_2192.n1 a_14262_2192.t4 5.8005
R3152 a_14262_2192.n1 a_14262_2192.t0 5.8005
R3153 a_14262_2192.n2 a_14262_2192.t2 5.8005
R3154 a_14262_2192.n2 a_14262_2192.t5 5.8005
R3155 a_14262_2192.n3 a_14262_2192.t7 5.8005
R3156 a_14262_2192.n3 a_14262_2192.t1 5.8005
R3157 a_14262_2192.n0 a_14262_2192.t9 5.8005
R3158 a_14262_2192.n0 a_14262_2192.t12 5.8005
R3159 a_14262_2192.n10 a_14262_2192.t8 5.8005
R3160 a_14262_2192.t11 a_14262_2192.n10 5.8005
R3161 a_14262_2192.n8 a_14262_2192.n6 1.94072
R3162 a_14262_2192.n9 a_14262_2192.n8 1.47876
R3163 a_14262_2192.n6 a_14262_2192.n5 0.478761
R3164 a_14262_2192.n5 a_14262_2192.n4 0.478761
R3165 a_2852_2192.n4 a_2852_2192.t12 32.0282
R3166 a_2852_2192.n10 a_2852_2192.n9 25.7663
R3167 a_2852_2192.n6 a_2852_2192.n1 25.75
R3168 a_2852_2192.n5 a_2852_2192.n2 25.75
R3169 a_2852_2192.n4 a_2852_2192.n3 25.75
R3170 a_2852_2192.n9 a_2852_2192.n0 25.288
R3171 a_2852_2192.n8 a_2852_2192.n7 24.288
R3172 a_2852_2192.n7 a_2852_2192.t4 5.8005
R3173 a_2852_2192.n7 a_2852_2192.t3 5.8005
R3174 a_2852_2192.n1 a_2852_2192.t1 5.8005
R3175 a_2852_2192.n1 a_2852_2192.t11 5.8005
R3176 a_2852_2192.n2 a_2852_2192.t9 5.8005
R3177 a_2852_2192.n2 a_2852_2192.t2 5.8005
R3178 a_2852_2192.n3 a_2852_2192.t0 5.8005
R3179 a_2852_2192.n3 a_2852_2192.t10 5.8005
R3180 a_2852_2192.n0 a_2852_2192.t7 5.8005
R3181 a_2852_2192.n0 a_2852_2192.t6 5.8005
R3182 a_2852_2192.t8 a_2852_2192.n10 5.8005
R3183 a_2852_2192.n10 a_2852_2192.t5 5.8005
R3184 a_2852_2192.n8 a_2852_2192.n6 1.94072
R3185 a_2852_2192.n9 a_2852_2192.n8 1.47876
R3186 a_2852_2192.n6 a_2852_2192.n5 0.478761
R3187 a_2852_2192.n5 a_2852_2192.n4 0.478761
R3188 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 879.481
R3189 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 742.783
R3190 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 665.16
R3191 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 623.388
R3192 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 523.774
R3193 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 431.807
R3194 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 427.875
R3195 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 357.26
R3196 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 208.537
R3197 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 168.077
R3198 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R3199 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R3200 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R3201 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 11.1806
R3202 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R3203 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R3204 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R3205 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R3206 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R3207 term_7.n1 term_7.t5 734.539
R3208 term_7.n1 term_7.t4 233.26
R3209 term_7.n2 term_7.n1 162.399
R3210 term_7.n2 term_7.n0 75.5108
R3211 term_7.n4 term_7.n3 66.3172
R3212 term_7.n3 term_7.t0 17.4005
R3213 term_7.n3 term_7.t2 17.4005
R3214 term_7.n0 term_7.t3 9.52217
R3215 term_7.n0 term_7.t1 9.52217
R3216 term_7 term_7.n4 5.08746
R3217 term_7.n4 term_7.n2 0.3755
R3218 saff_delay_unit_4/delay_unit_2_0.in_1.n1 saff_delay_unit_4/delay_unit_2_0.in_1.t14 572.12
R3219 saff_delay_unit_4/delay_unit_2_0.in_1.n1 saff_delay_unit_4/delay_unit_2_0.in_1.t9 572.12
R3220 saff_delay_unit_4/delay_unit_2_0.in_1.n0 saff_delay_unit_4/delay_unit_2_0.in_1.t16 572.12
R3221 saff_delay_unit_4/delay_unit_2_0.in_1.n0 saff_delay_unit_4/delay_unit_2_0.in_1.t10 572.12
R3222 saff_delay_unit_4/delay_unit_2_0.in_1.n6 saff_delay_unit_4/delay_unit_2_0.in_1.t13 523.774
R3223 saff_delay_unit_4/delay_unit_2_0.in_1.n7 saff_delay_unit_4/delay_unit_2_0.in_1.t18 523.774
R3224 saff_delay_unit_4/delay_unit_2_0.in_1.n3 saff_delay_unit_4/delay_unit_2_0.in_1.t17 523.774
R3225 saff_delay_unit_4/delay_unit_2_0.in_1.n4 saff_delay_unit_4/delay_unit_2_0.in_1.t19 523.774
R3226 saff_delay_unit_4/delay_unit_2_0.in_1.n6 saff_delay_unit_4/delay_unit_2_0.in_1.t15 202.44
R3227 saff_delay_unit_4/delay_unit_2_0.in_1.n7 saff_delay_unit_4/delay_unit_2_0.in_1.t11 202.44
R3228 saff_delay_unit_4/delay_unit_2_0.in_1.n3 saff_delay_unit_4/delay_unit_2_0.in_1.t8 202.44
R3229 saff_delay_unit_4/delay_unit_2_0.in_1.n4 saff_delay_unit_4/delay_unit_2_0.in_1.t12 202.44
R3230 saff_delay_unit_4/delay_unit_2_0.in_1.n2 saff_delay_unit_4/delay_unit_2_0.in_1.n0 166.468
R3231 saff_delay_unit_4/delay_unit_2_0.in_1.n9 saff_delay_unit_4/delay_unit_2_0.in_1.n5 166.149
R3232 saff_delay_unit_4/delay_unit_2_0.in_1.n9 saff_delay_unit_4/delay_unit_2_0.in_1.n8 165.8
R3233 saff_delay_unit_4/delay_unit_2_0.in_1.n2 saff_delay_unit_4/delay_unit_2_0.in_1.n1 165.8
R3234 saff_delay_unit_4/delay_unit_2_0.in_1.n10 saff_delay_unit_4/delay_unit_2_0.in_1.t6 85.1574
R3235 saff_delay_unit_4/delay_unit_2_0.in_1.n10 saff_delay_unit_4/delay_unit_2_0.in_1.t7 83.8097
R3236 saff_delay_unit_4/delay_unit_2_0.in_1.n16 saff_delay_unit_4/delay_unit_2_0.in_1.t5 83.8097
R3237 saff_delay_unit_4/delay_unit_2_0.in_1.n17 saff_delay_unit_4/delay_unit_2_0.in_1.t1 83.7172
R3238 saff_delay_unit_4/delay_unit_2_0.in_1.n14 saff_delay_unit_4/delay_unit_2_0.in_1.n13 74.288
R3239 saff_delay_unit_4/delay_unit_2_0.in_1.n14 saff_delay_unit_4/delay_unit_2_0.in_1.n12 67.7574
R3240 saff_delay_unit_4/delay_unit_2_0.in_1.n8 saff_delay_unit_4/delay_unit_2_0.in_1.n6 27.8082
R3241 saff_delay_unit_4/delay_unit_2_0.in_1.n5 saff_delay_unit_4/delay_unit_2_0.in_1.n4 27.8082
R3242 saff_delay_unit_4/delay_unit_2_0.in_1.n8 saff_delay_unit_4/delay_unit_2_0.in_1.n7 26.5723
R3243 saff_delay_unit_4/delay_unit_2_0.in_1.n5 saff_delay_unit_4/delay_unit_2_0.in_1.n3 26.5723
R3244 saff_delay_unit_4/delay_unit_2_0.in_1.n12 saff_delay_unit_4/delay_unit_2_0.in_1.t2 17.4005
R3245 saff_delay_unit_4/delay_unit_2_0.in_1.n12 saff_delay_unit_4/delay_unit_2_0.in_1.t0 17.4005
R3246 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_1.n2 16.0275
R3247 saff_delay_unit_4/delay_unit_2_0.in_1.n11 saff_delay_unit_4/delay_unit_2_0.in_1.n9 11.8364
R3248 saff_delay_unit_4/delay_unit_2_0.in_1.n13 saff_delay_unit_4/delay_unit_2_0.in_1.t3 9.52217
R3249 saff_delay_unit_4/delay_unit_2_0.in_1.n13 saff_delay_unit_4/delay_unit_2_0.in_1.t4 9.52217
R3250 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_1.n17 6.02878
R3251 saff_delay_unit_4/delay_unit_2_0.in_1.n15 saff_delay_unit_4/delay_unit_2_0.in_1.n14 5.83219
R3252 saff_delay_unit_4/delay_unit_2_0.in_1.n11 saff_delay_unit_4/delay_unit_2_0.in_1.n10 5.74235
R3253 saff_delay_unit_4/delay_unit_2_0.in_1.n16 saff_delay_unit_4/delay_unit_2_0.in_1.n15 5.49235
R3254 saff_delay_unit_4/delay_unit_2_0.in_1.n17 saff_delay_unit_4/delay_unit_2_0.in_1.n16 1.44072
R3255 saff_delay_unit_4/delay_unit_2_0.in_1.n15 saff_delay_unit_4/delay_unit_2_0.in_1 1.32081
R3256 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_1.n11 0.285656
R3257 saff_delay_unit_5/delay_unit_2_0.in_2.n8 saff_delay_unit_5/delay_unit_2_0.in_2.t8 784.053
R3258 saff_delay_unit_5/delay_unit_2_0.in_2.n8 saff_delay_unit_5/delay_unit_2_0.in_2.t13 784.053
R3259 saff_delay_unit_5/delay_unit_2_0.in_2.n9 saff_delay_unit_5/delay_unit_2_0.in_2.t12 784.053
R3260 saff_delay_unit_5/delay_unit_2_0.in_2.n9 saff_delay_unit_5/delay_unit_2_0.in_2.t17 784.053
R3261 saff_delay_unit_5/delay_unit_2_0.in_2.n3 saff_delay_unit_5/delay_unit_2_0.in_2.t16 523.774
R3262 saff_delay_unit_5/delay_unit_2_0.in_2.n4 saff_delay_unit_5/delay_unit_2_0.in_2.t10 523.774
R3263 saff_delay_unit_5/delay_unit_2_0.in_2.n0 saff_delay_unit_5/delay_unit_2_0.in_2.t18 523.774
R3264 saff_delay_unit_5/delay_unit_2_0.in_2.n1 saff_delay_unit_5/delay_unit_2_0.in_2.t11 523.774
R3265 saff_delay_unit_5/delay_unit_2_0.in_2.n3 saff_delay_unit_5/delay_unit_2_0.in_2.t19 202.44
R3266 saff_delay_unit_5/delay_unit_2_0.in_2.n4 saff_delay_unit_5/delay_unit_2_0.in_2.t14 202.44
R3267 saff_delay_unit_5/delay_unit_2_0.in_2.n0 saff_delay_unit_5/delay_unit_2_0.in_2.t9 202.44
R3268 saff_delay_unit_5/delay_unit_2_0.in_2.n1 saff_delay_unit_5/delay_unit_2_0.in_2.t15 202.44
R3269 saff_delay_unit_5/delay_unit_2_0.in_2.n10 saff_delay_unit_5/delay_unit_2_0.in_2.n8 168.659
R3270 saff_delay_unit_5/delay_unit_2_0.in_2.n10 saff_delay_unit_5/delay_unit_2_0.in_2.n9 167.992
R3271 saff_delay_unit_5/delay_unit_2_0.in_2.n6 saff_delay_unit_5/delay_unit_2_0.in_2.n2 166.144
R3272 saff_delay_unit_5/delay_unit_2_0.in_2.n6 saff_delay_unit_5/delay_unit_2_0.in_2.n5 165.8
R3273 saff_delay_unit_5/delay_unit_2_0.in_2.n14 saff_delay_unit_5/delay_unit_2_0.in_2.t4 85.2499
R3274 saff_delay_unit_5/delay_unit_2_0.in_2.n7 saff_delay_unit_5/delay_unit_2_0.in_2.t7 85.2499
R3275 saff_delay_unit_5/delay_unit_2_0.in_2.n14 saff_delay_unit_5/delay_unit_2_0.in_2.t2 83.7172
R3276 saff_delay_unit_5/delay_unit_2_0.in_2.n7 saff_delay_unit_5/delay_unit_2_0.in_2.t6 83.7172
R3277 saff_delay_unit_5/delay_unit_2_0.in_2.n13 saff_delay_unit_5/delay_unit_2_0.in_2.n11 75.7282
R3278 saff_delay_unit_5/delay_unit_2_0.in_2.n13 saff_delay_unit_5/delay_unit_2_0.in_2.n12 66.3172
R3279 saff_delay_unit_5/delay_unit_2_0.in_2.n5 saff_delay_unit_5/delay_unit_2_0.in_2.n3 27.8082
R3280 saff_delay_unit_5/delay_unit_2_0.in_2.n2 saff_delay_unit_5/delay_unit_2_0.in_2.n0 27.8082
R3281 saff_delay_unit_5/delay_unit_2_0.in_2.n5 saff_delay_unit_5/delay_unit_2_0.in_2.n4 26.5723
R3282 saff_delay_unit_5/delay_unit_2_0.in_2.n2 saff_delay_unit_5/delay_unit_2_0.in_2.n1 26.5723
R3283 saff_delay_unit_5/delay_unit_2_0.in_2.n12 saff_delay_unit_5/delay_unit_2_0.in_2.t1 17.4005
R3284 saff_delay_unit_5/delay_unit_2_0.in_2.n12 saff_delay_unit_5/delay_unit_2_0.in_2.t0 17.4005
R3285 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2.n10 17.1141
R3286 saff_delay_unit_5/delay_unit_2_0.in_2.n11 saff_delay_unit_5/delay_unit_2_0.in_2.t3 9.52217
R3287 saff_delay_unit_5/delay_unit_2_0.in_2.n11 saff_delay_unit_5/delay_unit_2_0.in_2.t5 9.52217
R3288 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2.n7 6.45821
R3289 saff_delay_unit_5/delay_unit_2_0.in_2.n15 saff_delay_unit_5/delay_unit_2_0.in_2.n13 5.30824
R3290 saff_delay_unit_5/delay_unit_2_0.in_2.n15 saff_delay_unit_5/delay_unit_2_0.in_2.n14 4.94887
R3291 saff_delay_unit_5/delay_unit_2_0.in_2.n16 saff_delay_unit_5/delay_unit_2_0.in_2 1.54347
R3292 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2.n6 1.06691
R3293 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2.n16 0.602062
R3294 saff_delay_unit_5/delay_unit_2_0.in_2.n16 saff_delay_unit_5/delay_unit_2_0.in_2 0.453625
R3295 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2.n15 0.160656
R3296 term_1.n1 term_1.t5 734.539
R3297 term_1.n1 term_1.t4 233.26
R3298 term_1.n2 term_1.n1 162.399
R3299 term_1.n2 term_1.n0 75.5108
R3300 term_1.n4 term_1.n3 66.3172
R3301 term_1.n3 term_1.t2 17.4005
R3302 term_1.n3 term_1.t0 17.4005
R3303 term_1.n0 term_1.t1 9.52217
R3304 term_1.n0 term_1.t3 9.52217
R3305 term_1 term_1.n4 5.08746
R3306 term_1.n4 term_1.n2 0.3755
R3307 saff_delay_unit_3/delay_unit_2_0.in_1.n12 saff_delay_unit_3/delay_unit_2_0.in_1.t12 572.12
R3308 saff_delay_unit_3/delay_unit_2_0.in_1.n12 saff_delay_unit_3/delay_unit_2_0.in_1.t18 572.12
R3309 saff_delay_unit_3/delay_unit_2_0.in_1.n11 saff_delay_unit_3/delay_unit_2_0.in_1.t14 572.12
R3310 saff_delay_unit_3/delay_unit_2_0.in_1.n11 saff_delay_unit_3/delay_unit_2_0.in_1.t19 572.12
R3311 saff_delay_unit_3/delay_unit_2_0.in_1.n3 saff_delay_unit_3/delay_unit_2_0.in_1.t8 523.774
R3312 saff_delay_unit_3/delay_unit_2_0.in_1.n4 saff_delay_unit_3/delay_unit_2_0.in_1.t13 523.774
R3313 saff_delay_unit_3/delay_unit_2_0.in_1.n0 saff_delay_unit_3/delay_unit_2_0.in_1.t9 523.774
R3314 saff_delay_unit_3/delay_unit_2_0.in_1.n1 saff_delay_unit_3/delay_unit_2_0.in_1.t15 523.774
R3315 saff_delay_unit_3/delay_unit_2_0.in_1.n3 saff_delay_unit_3/delay_unit_2_0.in_1.t10 202.44
R3316 saff_delay_unit_3/delay_unit_2_0.in_1.n4 saff_delay_unit_3/delay_unit_2_0.in_1.t16 202.44
R3317 saff_delay_unit_3/delay_unit_2_0.in_1.n0 saff_delay_unit_3/delay_unit_2_0.in_1.t11 202.44
R3318 saff_delay_unit_3/delay_unit_2_0.in_1.n1 saff_delay_unit_3/delay_unit_2_0.in_1.t17 202.44
R3319 saff_delay_unit_3/delay_unit_2_0.in_1.n13 saff_delay_unit_3/delay_unit_2_0.in_1.n11 166.468
R3320 saff_delay_unit_3/delay_unit_2_0.in_1.n6 saff_delay_unit_3/delay_unit_2_0.in_1.n2 166.149
R3321 saff_delay_unit_3/delay_unit_2_0.in_1.n13 saff_delay_unit_3/delay_unit_2_0.in_1.n12 165.8
R3322 saff_delay_unit_3/delay_unit_2_0.in_1.n6 saff_delay_unit_3/delay_unit_2_0.in_1.n5 165.8
R3323 saff_delay_unit_3/delay_unit_2_0.in_1.n7 saff_delay_unit_3/delay_unit_2_0.in_1.t6 85.1574
R3324 saff_delay_unit_3/delay_unit_2_0.in_1.n15 saff_delay_unit_3/delay_unit_2_0.in_1.t5 83.8097
R3325 saff_delay_unit_3/delay_unit_2_0.in_1.n7 saff_delay_unit_3/delay_unit_2_0.in_1.t7 83.8097
R3326 saff_delay_unit_3/delay_unit_2_0.in_1.n14 saff_delay_unit_3/delay_unit_2_0.in_1.t1 83.7172
R3327 saff_delay_unit_3/delay_unit_2_0.in_1.n10 saff_delay_unit_3/delay_unit_2_0.in_1.n9 74.288
R3328 saff_delay_unit_3/delay_unit_2_0.in_1.n10 saff_delay_unit_3/delay_unit_2_0.in_1.n8 67.7574
R3329 saff_delay_unit_3/delay_unit_2_0.in_1.n5 saff_delay_unit_3/delay_unit_2_0.in_1.n3 27.8082
R3330 saff_delay_unit_3/delay_unit_2_0.in_1.n2 saff_delay_unit_3/delay_unit_2_0.in_1.n1 27.8082
R3331 saff_delay_unit_3/delay_unit_2_0.in_1.n5 saff_delay_unit_3/delay_unit_2_0.in_1.n4 26.5723
R3332 saff_delay_unit_3/delay_unit_2_0.in_1.n2 saff_delay_unit_3/delay_unit_2_0.in_1.n0 26.5723
R3333 saff_delay_unit_3/delay_unit_2_0.in_1.n8 saff_delay_unit_3/delay_unit_2_0.in_1.t2 17.4005
R3334 saff_delay_unit_3/delay_unit_2_0.in_1.n8 saff_delay_unit_3/delay_unit_2_0.in_1.t4 17.4005
R3335 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_1.n13 16.0275
R3336 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_1.n6 11.8364
R3337 saff_delay_unit_3/delay_unit_2_0.in_1.n9 saff_delay_unit_3/delay_unit_2_0.in_1.t0 9.52217
R3338 saff_delay_unit_3/delay_unit_2_0.in_1.n9 saff_delay_unit_3/delay_unit_2_0.in_1.t3 9.52217
R3339 saff_delay_unit_3/delay_unit_2_0.in_1.n14 saff_delay_unit_3/delay_unit_2_0.in_1 6.02878
R3340 saff_delay_unit_3/delay_unit_2_0.in_1.n16 saff_delay_unit_3/delay_unit_2_0.in_1.n10 5.83219
R3341 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_1.n7 5.74235
R3342 saff_delay_unit_3/delay_unit_2_0.in_1.n16 saff_delay_unit_3/delay_unit_2_0.in_1.n15 5.49235
R3343 saff_delay_unit_3/delay_unit_2_0.in_1.n15 saff_delay_unit_3/delay_unit_2_0.in_1.n14 1.44072
R3344 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_1.n16 1.32081
R3345 a_16808_2192.n2 a_16808_2192.n1 34.9195
R3346 a_16808_2192.n3 a_16808_2192.n2 25.5407
R3347 a_16808_2192.n2 a_16808_2192.n0 25.2907
R3348 a_16808_2192.n1 a_16808_2192.t3 5.8005
R3349 a_16808_2192.n1 a_16808_2192.t1 5.8005
R3350 a_16808_2192.n0 a_16808_2192.t2 5.8005
R3351 a_16808_2192.n0 a_16808_2192.t0 5.8005
R3352 a_16808_2192.n3 a_16808_2192.t5 5.8005
R3353 a_16808_2192.t4 a_16808_2192.n3 5.8005
R3354 saff_delay_unit_2/delay_unit_2_0.in_2.n8 saff_delay_unit_2/delay_unit_2_0.in_2.t9 784.053
R3355 saff_delay_unit_2/delay_unit_2_0.in_2.n8 saff_delay_unit_2/delay_unit_2_0.in_2.t16 784.053
R3356 saff_delay_unit_2/delay_unit_2_0.in_2.n9 saff_delay_unit_2/delay_unit_2_0.in_2.t10 784.053
R3357 saff_delay_unit_2/delay_unit_2_0.in_2.n9 saff_delay_unit_2/delay_unit_2_0.in_2.t18 784.053
R3358 saff_delay_unit_2/delay_unit_2_0.in_2.n3 saff_delay_unit_2/delay_unit_2_0.in_2.t19 523.774
R3359 saff_delay_unit_2/delay_unit_2_0.in_2.n4 saff_delay_unit_2/delay_unit_2_0.in_2.t11 523.774
R3360 saff_delay_unit_2/delay_unit_2_0.in_2.n0 saff_delay_unit_2/delay_unit_2_0.in_2.t12 523.774
R3361 saff_delay_unit_2/delay_unit_2_0.in_2.n1 saff_delay_unit_2/delay_unit_2_0.in_2.t13 523.774
R3362 saff_delay_unit_2/delay_unit_2_0.in_2.n3 saff_delay_unit_2/delay_unit_2_0.in_2.t8 202.44
R3363 saff_delay_unit_2/delay_unit_2_0.in_2.n4 saff_delay_unit_2/delay_unit_2_0.in_2.t14 202.44
R3364 saff_delay_unit_2/delay_unit_2_0.in_2.n0 saff_delay_unit_2/delay_unit_2_0.in_2.t15 202.44
R3365 saff_delay_unit_2/delay_unit_2_0.in_2.n1 saff_delay_unit_2/delay_unit_2_0.in_2.t17 202.44
R3366 saff_delay_unit_2/delay_unit_2_0.in_2.n10 saff_delay_unit_2/delay_unit_2_0.in_2.n8 168.659
R3367 saff_delay_unit_2/delay_unit_2_0.in_2.n10 saff_delay_unit_2/delay_unit_2_0.in_2.n9 167.992
R3368 saff_delay_unit_2/delay_unit_2_0.in_2.n6 saff_delay_unit_2/delay_unit_2_0.in_2.n2 166.144
R3369 saff_delay_unit_2/delay_unit_2_0.in_2.n6 saff_delay_unit_2/delay_unit_2_0.in_2.n5 165.8
R3370 saff_delay_unit_2/delay_unit_2_0.in_2.n14 saff_delay_unit_2/delay_unit_2_0.in_2.t3 85.2499
R3371 saff_delay_unit_2/delay_unit_2_0.in_2.n7 saff_delay_unit_2/delay_unit_2_0.in_2.t7 85.2499
R3372 saff_delay_unit_2/delay_unit_2_0.in_2.n14 saff_delay_unit_2/delay_unit_2_0.in_2.t1 83.7172
R3373 saff_delay_unit_2/delay_unit_2_0.in_2.n7 saff_delay_unit_2/delay_unit_2_0.in_2.t6 83.7172
R3374 saff_delay_unit_2/delay_unit_2_0.in_2.n13 saff_delay_unit_2/delay_unit_2_0.in_2.n11 75.7282
R3375 saff_delay_unit_2/delay_unit_2_0.in_2.n13 saff_delay_unit_2/delay_unit_2_0.in_2.n12 66.3172
R3376 saff_delay_unit_2/delay_unit_2_0.in_2.n5 saff_delay_unit_2/delay_unit_2_0.in_2.n3 27.8082
R3377 saff_delay_unit_2/delay_unit_2_0.in_2.n2 saff_delay_unit_2/delay_unit_2_0.in_2.n0 27.8082
R3378 saff_delay_unit_2/delay_unit_2_0.in_2.n5 saff_delay_unit_2/delay_unit_2_0.in_2.n4 26.5723
R3379 saff_delay_unit_2/delay_unit_2_0.in_2.n2 saff_delay_unit_2/delay_unit_2_0.in_2.n1 26.5723
R3380 saff_delay_unit_2/delay_unit_2_0.in_2.n12 saff_delay_unit_2/delay_unit_2_0.in_2.t4 17.4005
R3381 saff_delay_unit_2/delay_unit_2_0.in_2.n12 saff_delay_unit_2/delay_unit_2_0.in_2.t0 17.4005
R3382 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n10 17.1141
R3383 saff_delay_unit_2/delay_unit_2_0.in_2.n11 saff_delay_unit_2/delay_unit_2_0.in_2.t5 9.52217
R3384 saff_delay_unit_2/delay_unit_2_0.in_2.n11 saff_delay_unit_2/delay_unit_2_0.in_2.t2 9.52217
R3385 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n7 6.45821
R3386 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n13 5.30824
R3387 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n14 4.94887
R3388 saff_delay_unit_2/delay_unit_2_0.in_2.n15 saff_delay_unit_2/delay_unit_2_0.in_2 1.70362
R3389 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n6 1.06691
R3390 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/delay_unit_2_0.in_2.n15 0.602062
R3391 saff_delay_unit_2/delay_unit_2_0.in_2.n15 saff_delay_unit_2/delay_unit_2_0.in_2 0.453625
R3392 saff_delay_unit_1/delay_unit_2_0.in_1.n13 saff_delay_unit_1/delay_unit_2_0.in_1.t15 572.12
R3393 saff_delay_unit_1/delay_unit_2_0.in_1.n13 saff_delay_unit_1/delay_unit_2_0.in_1.t8 572.12
R3394 saff_delay_unit_1/delay_unit_2_0.in_1.n12 saff_delay_unit_1/delay_unit_2_0.in_1.t18 572.12
R3395 saff_delay_unit_1/delay_unit_2_0.in_1.n12 saff_delay_unit_1/delay_unit_2_0.in_1.t14 572.12
R3396 saff_delay_unit_1/delay_unit_2_0.in_1.n3 saff_delay_unit_1/delay_unit_2_0.in_1.t16 523.774
R3397 saff_delay_unit_1/delay_unit_2_0.in_1.n4 saff_delay_unit_1/delay_unit_2_0.in_1.t9 523.774
R3398 saff_delay_unit_1/delay_unit_2_0.in_1.n0 saff_delay_unit_1/delay_unit_2_0.in_1.t13 523.774
R3399 saff_delay_unit_1/delay_unit_2_0.in_1.n1 saff_delay_unit_1/delay_unit_2_0.in_1.t10 523.774
R3400 saff_delay_unit_1/delay_unit_2_0.in_1.n3 saff_delay_unit_1/delay_unit_2_0.in_1.t19 202.44
R3401 saff_delay_unit_1/delay_unit_2_0.in_1.n4 saff_delay_unit_1/delay_unit_2_0.in_1.t11 202.44
R3402 saff_delay_unit_1/delay_unit_2_0.in_1.n0 saff_delay_unit_1/delay_unit_2_0.in_1.t17 202.44
R3403 saff_delay_unit_1/delay_unit_2_0.in_1.n1 saff_delay_unit_1/delay_unit_2_0.in_1.t12 202.44
R3404 saff_delay_unit_1/delay_unit_2_0.in_1.n14 saff_delay_unit_1/delay_unit_2_0.in_1.n12 166.468
R3405 saff_delay_unit_1/delay_unit_2_0.in_1.n6 saff_delay_unit_1/delay_unit_2_0.in_1.n2 166.149
R3406 saff_delay_unit_1/delay_unit_2_0.in_1.n14 saff_delay_unit_1/delay_unit_2_0.in_1.n13 165.8
R3407 saff_delay_unit_1/delay_unit_2_0.in_1.n6 saff_delay_unit_1/delay_unit_2_0.in_1.n5 165.8
R3408 saff_delay_unit_1/delay_unit_2_0.in_1.n7 saff_delay_unit_1/delay_unit_2_0.in_1.t6 85.1574
R3409 saff_delay_unit_1/delay_unit_2_0.in_1.n16 saff_delay_unit_1/delay_unit_2_0.in_1.t3 83.8097
R3410 saff_delay_unit_1/delay_unit_2_0.in_1.n7 saff_delay_unit_1/delay_unit_2_0.in_1.t7 83.8097
R3411 saff_delay_unit_1/delay_unit_2_0.in_1.n15 saff_delay_unit_1/delay_unit_2_0.in_1.t0 83.7172
R3412 saff_delay_unit_1/delay_unit_2_0.in_1.n11 saff_delay_unit_1/delay_unit_2_0.in_1.n10 74.288
R3413 saff_delay_unit_1/delay_unit_2_0.in_1.n11 saff_delay_unit_1/delay_unit_2_0.in_1.n9 67.7574
R3414 saff_delay_unit_1/delay_unit_2_0.in_1.n5 saff_delay_unit_1/delay_unit_2_0.in_1.n3 27.8082
R3415 saff_delay_unit_1/delay_unit_2_0.in_1.n2 saff_delay_unit_1/delay_unit_2_0.in_1.n1 27.8082
R3416 saff_delay_unit_1/delay_unit_2_0.in_1.n5 saff_delay_unit_1/delay_unit_2_0.in_1.n4 26.5723
R3417 saff_delay_unit_1/delay_unit_2_0.in_1.n2 saff_delay_unit_1/delay_unit_2_0.in_1.n0 26.5723
R3418 saff_delay_unit_1/delay_unit_2_0.in_1.n9 saff_delay_unit_1/delay_unit_2_0.in_1.t2 17.4005
R3419 saff_delay_unit_1/delay_unit_2_0.in_1.n9 saff_delay_unit_1/delay_unit_2_0.in_1.t1 17.4005
R3420 saff_delay_unit_1/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_1.n14 16.0275
R3421 saff_delay_unit_1/delay_unit_2_0.in_1.n8 saff_delay_unit_1/delay_unit_2_0.in_1.n6 11.8364
R3422 saff_delay_unit_1/delay_unit_2_0.in_1.n10 saff_delay_unit_1/delay_unit_2_0.in_1.t5 9.52217
R3423 saff_delay_unit_1/delay_unit_2_0.in_1.n10 saff_delay_unit_1/delay_unit_2_0.in_1.t4 9.52217
R3424 saff_delay_unit_1/delay_unit_2_0.in_1.n15 saff_delay_unit_1/delay_unit_2_0.in_1 6.02878
R3425 saff_delay_unit_1/delay_unit_2_0.in_1.n17 saff_delay_unit_1/delay_unit_2_0.in_1.n11 5.83219
R3426 saff_delay_unit_1/delay_unit_2_0.in_1.n8 saff_delay_unit_1/delay_unit_2_0.in_1.n7 5.74235
R3427 saff_delay_unit_1/delay_unit_2_0.in_1.n17 saff_delay_unit_1/delay_unit_2_0.in_1.n16 5.49235
R3428 saff_delay_unit_1/delay_unit_2_0.in_1.n16 saff_delay_unit_1/delay_unit_2_0.in_1.n15 1.44072
R3429 saff_delay_unit_1/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_1.n17 1.32081
R3430 saff_delay_unit_1/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_1.n8 0.285656
R3431 a_5134_2192.n6 a_5134_2192.t10 32.0282
R3432 a_5134_2192.n2 a_5134_2192.n1 25.7663
R3433 a_5134_2192.n8 a_5134_2192.n3 25.75
R3434 a_5134_2192.n7 a_5134_2192.n4 25.75
R3435 a_5134_2192.n6 a_5134_2192.n5 25.75
R3436 a_5134_2192.n2 a_5134_2192.n0 25.288
R3437 a_5134_2192.n10 a_5134_2192.n9 24.288
R3438 a_5134_2192.n0 a_5134_2192.t5 5.8005
R3439 a_5134_2192.n0 a_5134_2192.t4 5.8005
R3440 a_5134_2192.n1 a_5134_2192.t6 5.8005
R3441 a_5134_2192.n1 a_5134_2192.t7 5.8005
R3442 a_5134_2192.n3 a_5134_2192.t0 5.8005
R3443 a_5134_2192.n3 a_5134_2192.t11 5.8005
R3444 a_5134_2192.n4 a_5134_2192.t9 5.8005
R3445 a_5134_2192.n4 a_5134_2192.t3 5.8005
R3446 a_5134_2192.n5 a_5134_2192.t2 5.8005
R3447 a_5134_2192.n5 a_5134_2192.t12 5.8005
R3448 a_5134_2192.t8 a_5134_2192.n10 5.8005
R3449 a_5134_2192.n10 a_5134_2192.t1 5.8005
R3450 a_5134_2192.n9 a_5134_2192.n8 1.94072
R3451 a_5134_2192.n9 a_5134_2192.n2 1.47876
R3452 a_5134_2192.n8 a_5134_2192.n7 0.478761
R3453 a_5134_2192.n7 a_5134_2192.n6 0.478761
R3454 a_5398_2192.n2 a_5398_2192.n1 34.9195
R3455 a_5398_2192.n2 a_5398_2192.n0 25.5407
R3456 a_5398_2192.n3 a_5398_2192.n2 25.2907
R3457 a_5398_2192.n1 a_5398_2192.t3 5.8005
R3458 a_5398_2192.n1 a_5398_2192.t1 5.8005
R3459 a_5398_2192.n0 a_5398_2192.t5 5.8005
R3460 a_5398_2192.n0 a_5398_2192.t0 5.8005
R3461 a_5398_2192.n3 a_5398_2192.t2 5.8005
R3462 a_5398_2192.t4 a_5398_2192.n3 5.8005
R3463 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 879.481
R3464 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 742.783
R3465 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 665.16
R3466 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 623.388
R3467 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 523.774
R3468 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 431.807
R3469 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 427.875
R3470 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 357.26
R3471 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 208.537
R3472 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 168.077
R3473 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R3474 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R3475 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 31.2347
R3476 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 11.1806
R3477 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R3478 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R3479 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R3480 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R3481 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R3482 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 890.727
R3483 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 742.783
R3484 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 665.16
R3485 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 623.388
R3486 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 523.774
R3487 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 431.807
R3488 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 427.875
R3489 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 364.733
R3490 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 208.5
R3491 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 168.007
R3492 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R3493 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 31.2728
R3494 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 31.0337
R3495 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3496 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R3497 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 9.08234
R3498 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R3499 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R3500 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3501 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R3502 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R3503 saff_delay_unit_7/delay_unit_2_0.in_2.n8 saff_delay_unit_7/delay_unit_2_0.in_2.t17 784.053
R3504 saff_delay_unit_7/delay_unit_2_0.in_2.n8 saff_delay_unit_7/delay_unit_2_0.in_2.t10 784.053
R3505 saff_delay_unit_7/delay_unit_2_0.in_2.n9 saff_delay_unit_7/delay_unit_2_0.in_2.t18 784.053
R3506 saff_delay_unit_7/delay_unit_2_0.in_2.n9 saff_delay_unit_7/delay_unit_2_0.in_2.t11 784.053
R3507 saff_delay_unit_7/delay_unit_2_0.in_2.n3 saff_delay_unit_7/delay_unit_2_0.in_2.t14 523.774
R3508 saff_delay_unit_7/delay_unit_2_0.in_2.n4 saff_delay_unit_7/delay_unit_2_0.in_2.t9 523.774
R3509 saff_delay_unit_7/delay_unit_2_0.in_2.n0 saff_delay_unit_7/delay_unit_2_0.in_2.t19 523.774
R3510 saff_delay_unit_7/delay_unit_2_0.in_2.n1 saff_delay_unit_7/delay_unit_2_0.in_2.t12 523.774
R3511 saff_delay_unit_7/delay_unit_2_0.in_2.n3 saff_delay_unit_7/delay_unit_2_0.in_2.t16 202.44
R3512 saff_delay_unit_7/delay_unit_2_0.in_2.n4 saff_delay_unit_7/delay_unit_2_0.in_2.t13 202.44
R3513 saff_delay_unit_7/delay_unit_2_0.in_2.n0 saff_delay_unit_7/delay_unit_2_0.in_2.t8 202.44
R3514 saff_delay_unit_7/delay_unit_2_0.in_2.n1 saff_delay_unit_7/delay_unit_2_0.in_2.t15 202.44
R3515 saff_delay_unit_7/delay_unit_2_0.in_2.n10 saff_delay_unit_7/delay_unit_2_0.in_2.n8 168.659
R3516 saff_delay_unit_7/delay_unit_2_0.in_2.n10 saff_delay_unit_7/delay_unit_2_0.in_2.n9 167.992
R3517 saff_delay_unit_7/delay_unit_2_0.in_2.n6 saff_delay_unit_7/delay_unit_2_0.in_2.n2 166.144
R3518 saff_delay_unit_7/delay_unit_2_0.in_2.n6 saff_delay_unit_7/delay_unit_2_0.in_2.n5 165.8
R3519 saff_delay_unit_7/delay_unit_2_0.in_2.n14 saff_delay_unit_7/delay_unit_2_0.in_2.t5 85.2499
R3520 saff_delay_unit_7/delay_unit_2_0.in_2.n7 saff_delay_unit_7/delay_unit_2_0.in_2.t2 85.2499
R3521 saff_delay_unit_7/delay_unit_2_0.in_2.n7 saff_delay_unit_7/delay_unit_2_0.in_2.t1 83.7172
R3522 saff_delay_unit_7/delay_unit_2_0.in_2.n14 saff_delay_unit_7/delay_unit_2_0.in_2.t0 83.7172
R3523 saff_delay_unit_7/delay_unit_2_0.in_2.n13 saff_delay_unit_7/delay_unit_2_0.in_2.n11 75.7282
R3524 saff_delay_unit_7/delay_unit_2_0.in_2.n13 saff_delay_unit_7/delay_unit_2_0.in_2.n12 66.3172
R3525 saff_delay_unit_7/delay_unit_2_0.in_2.n5 saff_delay_unit_7/delay_unit_2_0.in_2.n3 27.8082
R3526 saff_delay_unit_7/delay_unit_2_0.in_2.n2 saff_delay_unit_7/delay_unit_2_0.in_2.n0 27.8082
R3527 saff_delay_unit_7/delay_unit_2_0.in_2.n5 saff_delay_unit_7/delay_unit_2_0.in_2.n4 26.5723
R3528 saff_delay_unit_7/delay_unit_2_0.in_2.n2 saff_delay_unit_7/delay_unit_2_0.in_2.n1 26.5723
R3529 saff_delay_unit_7/delay_unit_2_0.in_2.n12 saff_delay_unit_7/delay_unit_2_0.in_2.t7 17.4005
R3530 saff_delay_unit_7/delay_unit_2_0.in_2.n12 saff_delay_unit_7/delay_unit_2_0.in_2.t3 17.4005
R3531 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n10 17.1141
R3532 saff_delay_unit_7/delay_unit_2_0.in_2.n11 saff_delay_unit_7/delay_unit_2_0.in_2.t4 9.52217
R3533 saff_delay_unit_7/delay_unit_2_0.in_2.n11 saff_delay_unit_7/delay_unit_2_0.in_2.t6 9.52217
R3534 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n7 6.45821
R3535 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n13 5.30824
R3536 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n14 4.94887
R3537 saff_delay_unit_7/delay_unit_2_0.in_2.n15 saff_delay_unit_7/delay_unit_2_0.in_2 1.70362
R3538 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n6 1.06691
R3539 saff_delay_unit_7/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2.n15 0.602062
R3540 saff_delay_unit_7/delay_unit_2_0.in_2.n15 saff_delay_unit_7/delay_unit_2_0.in_2 0.453625
R3541 term_5.n1 term_5.t5 734.539
R3542 term_5.n1 term_5.t4 233.26
R3543 term_5.n2 term_5.n1 162.399
R3544 term_5.n2 term_5.n0 75.5108
R3545 term_5.n4 term_5.n3 66.3172
R3546 term_5.n3 term_5.t3 17.4005
R3547 term_5.n3 term_5.t1 17.4005
R3548 term_5.n0 term_5.t2 9.52217
R3549 term_5.n0 term_5.t0 9.52217
R3550 term_5 term_5.n4 5.08746
R3551 term_5.n4 term_5.n2 0.3755
R3552 saff_delay_unit_6/delay_unit_2_0.in_2.n8 saff_delay_unit_6/delay_unit_2_0.in_2.t10 784.053
R3553 saff_delay_unit_6/delay_unit_2_0.in_2.n8 saff_delay_unit_6/delay_unit_2_0.in_2.t17 784.053
R3554 saff_delay_unit_6/delay_unit_2_0.in_2.n9 saff_delay_unit_6/delay_unit_2_0.in_2.t14 784.053
R3555 saff_delay_unit_6/delay_unit_2_0.in_2.n9 saff_delay_unit_6/delay_unit_2_0.in_2.t19 784.053
R3556 saff_delay_unit_6/delay_unit_2_0.in_2.n3 saff_delay_unit_6/delay_unit_2_0.in_2.t9 523.774
R3557 saff_delay_unit_6/delay_unit_2_0.in_2.n4 saff_delay_unit_6/delay_unit_2_0.in_2.t11 523.774
R3558 saff_delay_unit_6/delay_unit_2_0.in_2.n0 saff_delay_unit_6/delay_unit_2_0.in_2.t12 523.774
R3559 saff_delay_unit_6/delay_unit_2_0.in_2.n1 saff_delay_unit_6/delay_unit_2_0.in_2.t18 523.774
R3560 saff_delay_unit_6/delay_unit_2_0.in_2.n3 saff_delay_unit_6/delay_unit_2_0.in_2.t13 202.44
R3561 saff_delay_unit_6/delay_unit_2_0.in_2.n4 saff_delay_unit_6/delay_unit_2_0.in_2.t15 202.44
R3562 saff_delay_unit_6/delay_unit_2_0.in_2.n0 saff_delay_unit_6/delay_unit_2_0.in_2.t16 202.44
R3563 saff_delay_unit_6/delay_unit_2_0.in_2.n1 saff_delay_unit_6/delay_unit_2_0.in_2.t8 202.44
R3564 saff_delay_unit_6/delay_unit_2_0.in_2.n10 saff_delay_unit_6/delay_unit_2_0.in_2.n8 168.659
R3565 saff_delay_unit_6/delay_unit_2_0.in_2.n10 saff_delay_unit_6/delay_unit_2_0.in_2.n9 167.992
R3566 saff_delay_unit_6/delay_unit_2_0.in_2.n6 saff_delay_unit_6/delay_unit_2_0.in_2.n2 166.144
R3567 saff_delay_unit_6/delay_unit_2_0.in_2.n6 saff_delay_unit_6/delay_unit_2_0.in_2.n5 165.8
R3568 saff_delay_unit_6/delay_unit_2_0.in_2.n14 saff_delay_unit_6/delay_unit_2_0.in_2.t4 85.2499
R3569 saff_delay_unit_6/delay_unit_2_0.in_2.n7 saff_delay_unit_6/delay_unit_2_0.in_2.t7 85.2499
R3570 saff_delay_unit_6/delay_unit_2_0.in_2.n14 saff_delay_unit_6/delay_unit_2_0.in_2.t2 83.7172
R3571 saff_delay_unit_6/delay_unit_2_0.in_2.n7 saff_delay_unit_6/delay_unit_2_0.in_2.t0 83.7172
R3572 saff_delay_unit_6/delay_unit_2_0.in_2.n13 saff_delay_unit_6/delay_unit_2_0.in_2.n11 75.7282
R3573 saff_delay_unit_6/delay_unit_2_0.in_2.n13 saff_delay_unit_6/delay_unit_2_0.in_2.n12 66.3172
R3574 saff_delay_unit_6/delay_unit_2_0.in_2.n5 saff_delay_unit_6/delay_unit_2_0.in_2.n3 27.8082
R3575 saff_delay_unit_6/delay_unit_2_0.in_2.n2 saff_delay_unit_6/delay_unit_2_0.in_2.n0 27.8082
R3576 saff_delay_unit_6/delay_unit_2_0.in_2.n5 saff_delay_unit_6/delay_unit_2_0.in_2.n4 26.5723
R3577 saff_delay_unit_6/delay_unit_2_0.in_2.n2 saff_delay_unit_6/delay_unit_2_0.in_2.n1 26.5723
R3578 saff_delay_unit_6/delay_unit_2_0.in_2.n12 saff_delay_unit_6/delay_unit_2_0.in_2.t1 17.4005
R3579 saff_delay_unit_6/delay_unit_2_0.in_2.n12 saff_delay_unit_6/delay_unit_2_0.in_2.t3 17.4005
R3580 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/delay_unit_2_0.in_2.n10 17.1141
R3581 saff_delay_unit_6/delay_unit_2_0.in_2.n11 saff_delay_unit_6/delay_unit_2_0.in_2.t6 9.52217
R3582 saff_delay_unit_6/delay_unit_2_0.in_2.n11 saff_delay_unit_6/delay_unit_2_0.in_2.t5 9.52217
R3583 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/delay_unit_2_0.in_2.n7 6.45821
R3584 saff_delay_unit_6/delay_unit_2_0.in_2.n15 saff_delay_unit_6/delay_unit_2_0.in_2.n13 5.30824
R3585 saff_delay_unit_6/delay_unit_2_0.in_2.n15 saff_delay_unit_6/delay_unit_2_0.in_2.n14 4.94887
R3586 saff_delay_unit_6/delay_unit_2_0.in_2.n16 saff_delay_unit_6/delay_unit_2_0.in_2 1.54347
R3587 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/delay_unit_2_0.in_2.n6 1.06691
R3588 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/delay_unit_2_0.in_2.n16 0.602062
R3589 saff_delay_unit_6/delay_unit_2_0.in_2.n16 saff_delay_unit_6/delay_unit_2_0.in_2 0.453625
R3590 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/delay_unit_2_0.in_2.n15 0.160656
R3591 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 890.727
R3592 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 742.783
R3593 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 665.16
R3594 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 623.388
R3595 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 523.774
R3596 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 431.807
R3597 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 427.875
R3598 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 364.733
R3599 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 208.5
R3600 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 168.007
R3601 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 75.2663
R3602 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 31.2728
R3603 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R3604 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3605 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R3606 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 9.08234
R3607 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R3608 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 4.50239
R3609 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 0.898227
R3610 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 0.707022
R3611 a_7416_2192.n4 a_7416_2192.t3 32.0282
R3612 a_7416_2192.n9 a_7416_2192.n0 25.7663
R3613 a_7416_2192.n6 a_7416_2192.n1 25.75
R3614 a_7416_2192.n5 a_7416_2192.n2 25.75
R3615 a_7416_2192.n4 a_7416_2192.n3 25.75
R3616 a_7416_2192.n10 a_7416_2192.n9 25.288
R3617 a_7416_2192.n8 a_7416_2192.n7 24.288
R3618 a_7416_2192.n7 a_7416_2192.t6 5.8005
R3619 a_7416_2192.n7 a_7416_2192.t9 5.8005
R3620 a_7416_2192.n1 a_7416_2192.t10 5.8005
R3621 a_7416_2192.n1 a_7416_2192.t0 5.8005
R3622 a_7416_2192.n2 a_7416_2192.t2 5.8005
R3623 a_7416_2192.n2 a_7416_2192.t11 5.8005
R3624 a_7416_2192.n3 a_7416_2192.t12 5.8005
R3625 a_7416_2192.n3 a_7416_2192.t1 5.8005
R3626 a_7416_2192.n0 a_7416_2192.t4 5.8005
R3627 a_7416_2192.n0 a_7416_2192.t7 5.8005
R3628 a_7416_2192.n10 a_7416_2192.t5 5.8005
R3629 a_7416_2192.t8 a_7416_2192.n10 5.8005
R3630 a_7416_2192.n8 a_7416_2192.n6 1.94072
R3631 a_7416_2192.n9 a_7416_2192.n8 1.47876
R3632 a_7416_2192.n6 a_7416_2192.n5 0.478761
R3633 a_7416_2192.n5 a_7416_2192.n4 0.478761
R3634 saff_delay_unit_7/saff_2_0.nd.n0 saff_delay_unit_7/saff_2_0.nd.t17 784.053
R3635 saff_delay_unit_7/saff_2_0.nd.n0 saff_delay_unit_7/saff_2_0.nd.t12 784.053
R3636 saff_delay_unit_7/saff_2_0.nd.n1 saff_delay_unit_7/saff_2_0.nd.t10 784.053
R3637 saff_delay_unit_7/saff_2_0.nd.n1 saff_delay_unit_7/saff_2_0.nd.t18 784.053
R3638 saff_delay_unit_7/saff_2_0.nd.n6 saff_delay_unit_7/saff_2_0.nd.t8 523.774
R3639 saff_delay_unit_7/saff_2_0.nd.n7 saff_delay_unit_7/saff_2_0.nd.t11 523.774
R3640 saff_delay_unit_7/saff_2_0.nd.n3 saff_delay_unit_7/saff_2_0.nd.t19 523.774
R3641 saff_delay_unit_7/saff_2_0.nd.n4 saff_delay_unit_7/saff_2_0.nd.t14 523.774
R3642 saff_delay_unit_7/saff_2_0.nd.n6 saff_delay_unit_7/saff_2_0.nd.t13 202.44
R3643 saff_delay_unit_7/saff_2_0.nd.n7 saff_delay_unit_7/saff_2_0.nd.t15 202.44
R3644 saff_delay_unit_7/saff_2_0.nd.n3 saff_delay_unit_7/saff_2_0.nd.t9 202.44
R3645 saff_delay_unit_7/saff_2_0.nd.n4 saff_delay_unit_7/saff_2_0.nd.t16 202.44
R3646 saff_delay_unit_7/saff_2_0.nd.n2 saff_delay_unit_7/saff_2_0.nd.n0 168.659
R3647 saff_delay_unit_7/saff_2_0.nd.n2 saff_delay_unit_7/saff_2_0.nd.n1 167.992
R3648 saff_delay_unit_7/saff_2_0.nd.n9 saff_delay_unit_7/saff_2_0.nd.n5 166.144
R3649 saff_delay_unit_7/saff_2_0.nd.n9 saff_delay_unit_7/saff_2_0.nd.n8 165.8
R3650 saff_delay_unit_7/saff_2_0.nd.n15 saff_delay_unit_7/saff_2_0.nd.t4 85.2499
R3651 saff_delay_unit_7/saff_2_0.nd.n10 saff_delay_unit_7/saff_2_0.nd.t7 85.2499
R3652 saff_delay_unit_7/saff_2_0.nd.n15 saff_delay_unit_7/saff_2_0.nd.t2 83.7172
R3653 saff_delay_unit_7/saff_2_0.nd.n10 saff_delay_unit_7/saff_2_0.nd.t6 83.7172
R3654 saff_delay_unit_7/saff_2_0.nd.n14 saff_delay_unit_7/saff_2_0.nd.n12 75.7282
R3655 saff_delay_unit_7/saff_2_0.nd.n14 saff_delay_unit_7/saff_2_0.nd.n13 66.3172
R3656 saff_delay_unit_7/saff_2_0.nd.n8 saff_delay_unit_7/saff_2_0.nd.n6 27.8082
R3657 saff_delay_unit_7/saff_2_0.nd.n5 saff_delay_unit_7/saff_2_0.nd.n3 27.8082
R3658 saff_delay_unit_7/saff_2_0.nd.n8 saff_delay_unit_7/saff_2_0.nd.n7 26.5723
R3659 saff_delay_unit_7/saff_2_0.nd.n5 saff_delay_unit_7/saff_2_0.nd.n4 26.5723
R3660 saff_delay_unit_7/saff_2_0.nd.n13 saff_delay_unit_7/saff_2_0.nd.t1 17.4005
R3661 saff_delay_unit_7/saff_2_0.nd.n13 saff_delay_unit_7/saff_2_0.nd.t0 17.4005
R3662 saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd saff_delay_unit_7/saff_2_0.nd.n2 17.1141
R3663 saff_delay_unit_7/saff_2_0.nd.n12 saff_delay_unit_7/saff_2_0.nd.t3 9.52217
R3664 saff_delay_unit_7/saff_2_0.nd.n12 saff_delay_unit_7/saff_2_0.nd.t5 9.52217
R3665 delay_unit_2_0.in_2 saff_delay_unit_7/saff_2_0.nd.n10 6.45821
R3666 saff_delay_unit_7/saff_2_0.nd.n16 saff_delay_unit_7/saff_2_0.nd.n14 5.30824
R3667 saff_delay_unit_7/saff_2_0.nd.n16 saff_delay_unit_7/saff_2_0.nd.n15 4.94887
R3668 saff_delay_unit_7/delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.nd.n11 1.54347
R3669 delay_unit_2_0.in_2 saff_delay_unit_7/saff_2_0.nd.n9 1.06691
R3670 saff_delay_unit_7/saff_2_0.nd.n11 delay_unit_2_0.in_2 0.602062
R3671 saff_delay_unit_7/saff_2_0.nd.n11 saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd 0.453625
R3672 saff_delay_unit_7/delay_unit_2_0.out_2 saff_delay_unit_7/saff_2_0.nd.n16 0.160656
R3673 delay_unit_2_0.out_1.n3 delay_unit_2_0.out_1.t2 85.1574
R3674 delay_unit_2_0.out_1.n3 delay_unit_2_0.out_1.t3 83.8097
R3675 delay_unit_2_0.out_1.n2 delay_unit_2_0.out_1.n1 74.288
R3676 delay_unit_2_0.out_1.n2 delay_unit_2_0.out_1.n0 67.7574
R3677 delay_unit_2_0.out_1.n0 delay_unit_2_0.out_1.t0 17.4005
R3678 delay_unit_2_0.out_1.n0 delay_unit_2_0.out_1.t1 17.4005
R3679 delay_unit_2_0.out_1.n1 delay_unit_2_0.out_1.t4 9.52217
R3680 delay_unit_2_0.out_1.n1 delay_unit_2_0.out_1.t5 9.52217
R3681 delay_unit_2_0.out_1.n4 delay_unit_2_0.out_1.n2 5.83219
R3682 delay_unit_2_0.out_1.n4 delay_unit_2_0.out_1.n3 5.49235
R3683 delay_unit_2_0.out_1 delay_unit_2_0.out_1.n4 1.32081
R3684 saff_delay_unit_6/delay_unit_2_0.in_1.n13 saff_delay_unit_6/delay_unit_2_0.in_1.t11 572.12
R3685 saff_delay_unit_6/delay_unit_2_0.in_1.n13 saff_delay_unit_6/delay_unit_2_0.in_1.t16 572.12
R3686 saff_delay_unit_6/delay_unit_2_0.in_1.n12 saff_delay_unit_6/delay_unit_2_0.in_1.t14 572.12
R3687 saff_delay_unit_6/delay_unit_2_0.in_1.n12 saff_delay_unit_6/delay_unit_2_0.in_1.t9 572.12
R3688 saff_delay_unit_6/delay_unit_2_0.in_1.n3 saff_delay_unit_6/delay_unit_2_0.in_1.t12 523.774
R3689 saff_delay_unit_6/delay_unit_2_0.in_1.n4 saff_delay_unit_6/delay_unit_2_0.in_1.t17 523.774
R3690 saff_delay_unit_6/delay_unit_2_0.in_1.n0 saff_delay_unit_6/delay_unit_2_0.in_1.t10 523.774
R3691 saff_delay_unit_6/delay_unit_2_0.in_1.n1 saff_delay_unit_6/delay_unit_2_0.in_1.t18 523.774
R3692 saff_delay_unit_6/delay_unit_2_0.in_1.n3 saff_delay_unit_6/delay_unit_2_0.in_1.t15 202.44
R3693 saff_delay_unit_6/delay_unit_2_0.in_1.n4 saff_delay_unit_6/delay_unit_2_0.in_1.t19 202.44
R3694 saff_delay_unit_6/delay_unit_2_0.in_1.n0 saff_delay_unit_6/delay_unit_2_0.in_1.t13 202.44
R3695 saff_delay_unit_6/delay_unit_2_0.in_1.n1 saff_delay_unit_6/delay_unit_2_0.in_1.t8 202.44
R3696 saff_delay_unit_6/delay_unit_2_0.in_1.n14 saff_delay_unit_6/delay_unit_2_0.in_1.n12 166.468
R3697 saff_delay_unit_6/delay_unit_2_0.in_1.n6 saff_delay_unit_6/delay_unit_2_0.in_1.n2 166.149
R3698 saff_delay_unit_6/delay_unit_2_0.in_1.n14 saff_delay_unit_6/delay_unit_2_0.in_1.n13 165.8
R3699 saff_delay_unit_6/delay_unit_2_0.in_1.n6 saff_delay_unit_6/delay_unit_2_0.in_1.n5 165.8
R3700 saff_delay_unit_6/delay_unit_2_0.in_1.n7 saff_delay_unit_6/delay_unit_2_0.in_1.t0 85.1574
R3701 saff_delay_unit_6/delay_unit_2_0.in_1.n16 saff_delay_unit_6/delay_unit_2_0.in_1.t5 83.8097
R3702 saff_delay_unit_6/delay_unit_2_0.in_1.n7 saff_delay_unit_6/delay_unit_2_0.in_1.t1 83.8097
R3703 saff_delay_unit_6/delay_unit_2_0.in_1.n15 saff_delay_unit_6/delay_unit_2_0.in_1.t4 83.7172
R3704 saff_delay_unit_6/delay_unit_2_0.in_1.n11 saff_delay_unit_6/delay_unit_2_0.in_1.n10 74.288
R3705 saff_delay_unit_6/delay_unit_2_0.in_1.n11 saff_delay_unit_6/delay_unit_2_0.in_1.n9 67.7574
R3706 saff_delay_unit_6/delay_unit_2_0.in_1.n5 saff_delay_unit_6/delay_unit_2_0.in_1.n3 27.8082
R3707 saff_delay_unit_6/delay_unit_2_0.in_1.n2 saff_delay_unit_6/delay_unit_2_0.in_1.n1 27.8082
R3708 saff_delay_unit_6/delay_unit_2_0.in_1.n5 saff_delay_unit_6/delay_unit_2_0.in_1.n4 26.5723
R3709 saff_delay_unit_6/delay_unit_2_0.in_1.n2 saff_delay_unit_6/delay_unit_2_0.in_1.n0 26.5723
R3710 saff_delay_unit_6/delay_unit_2_0.in_1.n9 saff_delay_unit_6/delay_unit_2_0.in_1.t3 17.4005
R3711 saff_delay_unit_6/delay_unit_2_0.in_1.n9 saff_delay_unit_6/delay_unit_2_0.in_1.t2 17.4005
R3712 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_6/delay_unit_2_0.in_1.n14 16.0275
R3713 saff_delay_unit_6/delay_unit_2_0.in_1.n8 saff_delay_unit_6/delay_unit_2_0.in_1.n6 11.8364
R3714 saff_delay_unit_6/delay_unit_2_0.in_1.n10 saff_delay_unit_6/delay_unit_2_0.in_1.t7 9.52217
R3715 saff_delay_unit_6/delay_unit_2_0.in_1.n10 saff_delay_unit_6/delay_unit_2_0.in_1.t6 9.52217
R3716 saff_delay_unit_6/delay_unit_2_0.in_1.n15 saff_delay_unit_6/delay_unit_2_0.in_1 6.02878
R3717 saff_delay_unit_6/delay_unit_2_0.in_1.n17 saff_delay_unit_6/delay_unit_2_0.in_1.n11 5.83219
R3718 saff_delay_unit_6/delay_unit_2_0.in_1.n8 saff_delay_unit_6/delay_unit_2_0.in_1.n7 5.74235
R3719 saff_delay_unit_6/delay_unit_2_0.in_1.n17 saff_delay_unit_6/delay_unit_2_0.in_1.n16 5.49235
R3720 saff_delay_unit_6/delay_unit_2_0.in_1.n16 saff_delay_unit_6/delay_unit_2_0.in_1.n15 1.44072
R3721 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_6/delay_unit_2_0.in_1.n17 1.32081
R3722 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_6/delay_unit_2_0.in_1.n8 0.285656
R3723 a_9962_2192.n2 a_9962_2192.n1 34.9195
R3724 a_9962_2192.n3 a_9962_2192.n2 25.5407
R3725 a_9962_2192.n2 a_9962_2192.n0 25.2907
R3726 a_9962_2192.n1 a_9962_2192.t0 5.8005
R3727 a_9962_2192.n1 a_9962_2192.t1 5.8005
R3728 a_9962_2192.n0 a_9962_2192.t2 5.8005
R3729 a_9962_2192.n0 a_9962_2192.t3 5.8005
R3730 a_9962_2192.n3 a_9962_2192.t5 5.8005
R3731 a_9962_2192.t4 a_9962_2192.n3 5.8005
R3732 a_9698_2192.n4 a_9698_2192.t2 32.0282
R3733 a_9698_2192.n9 a_9698_2192.n0 25.7663
R3734 a_9698_2192.n6 a_9698_2192.n1 25.75
R3735 a_9698_2192.n5 a_9698_2192.n2 25.75
R3736 a_9698_2192.n4 a_9698_2192.n3 25.75
R3737 a_9698_2192.n10 a_9698_2192.n9 25.288
R3738 a_9698_2192.n8 a_9698_2192.n7 24.288
R3739 a_9698_2192.n7 a_9698_2192.t5 5.8005
R3740 a_9698_2192.n7 a_9698_2192.t11 5.8005
R3741 a_9698_2192.n1 a_9698_2192.t9 5.8005
R3742 a_9698_2192.n1 a_9698_2192.t3 5.8005
R3743 a_9698_2192.n2 a_9698_2192.t1 5.8005
R3744 a_9698_2192.n2 a_9698_2192.t12 5.8005
R3745 a_9698_2192.n3 a_9698_2192.t10 5.8005
R3746 a_9698_2192.n3 a_9698_2192.t0 5.8005
R3747 a_9698_2192.n0 a_9698_2192.t4 5.8005
R3748 a_9698_2192.n0 a_9698_2192.t7 5.8005
R3749 a_9698_2192.n10 a_9698_2192.t6 5.8005
R3750 a_9698_2192.t8 a_9698_2192.n10 5.8005
R3751 a_9698_2192.n8 a_9698_2192.n6 1.94072
R3752 a_9698_2192.n9 a_9698_2192.n8 1.47876
R3753 a_9698_2192.n6 a_9698_2192.n5 0.478761
R3754 a_9698_2192.n5 a_9698_2192.n4 0.478761
R3755 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 879.481
R3756 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 742.783
R3757 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 665.16
R3758 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 623.388
R3759 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 523.774
R3760 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 431.807
R3761 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 427.875
R3762 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 357.26
R3763 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 208.537
R3764 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 168.077
R3765 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 75.5326
R3766 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R3767 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R3768 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 11.1806
R3769 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 10.5958
R3770 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R3771 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R3772 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 0.803118
R3773 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 0.23963
R3774 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 0.23963
R3775 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 890.727
R3776 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 742.783
R3777 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 665.16
R3778 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 623.388
R3779 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 523.774
R3780 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 431.807
R3781 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 427.875
R3782 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 364.733
R3783 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 208.5
R3784 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 168.007
R3785 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R3786 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 31.2728
R3787 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R3788 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R3789 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R3790 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R3791 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 8.00471
R3792 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R3793 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3794 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R3795 term_0.n1 term_0.t5 734.539
R3796 term_0.n1 term_0.t4 233.26
R3797 term_0.n2 term_0.n1 162.399
R3798 term_0.n2 term_0.n0 75.5108
R3799 term_0.n4 term_0.n3 66.3172
R3800 term_0.n3 term_0.t0 17.4005
R3801 term_0.n3 term_0.t1 17.4005
R3802 term_0.n0 term_0.t2 9.52217
R3803 term_0.n0 term_0.t3 9.52217
R3804 term_0 term_0.n4 5.08746
R3805 term_0.n4 term_0.n2 0.3755
R3806 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 890.727
R3807 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 742.783
R3808 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 665.16
R3809 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 623.388
R3810 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 523.774
R3811 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 431.807
R3812 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 427.875
R3813 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 364.733
R3814 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 208.5
R3815 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 168.007
R3816 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R3817 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 31.2728
R3818 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R3819 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R3820 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3821 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 9.08234
R3822 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R3823 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R3824 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3825 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R3826 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R3827 a_14526_2192.n2 a_14526_2192.n1 34.9195
R3828 a_14526_2192.n2 a_14526_2192.n0 25.5407
R3829 a_14526_2192.n3 a_14526_2192.n2 25.2907
R3830 a_14526_2192.n1 a_14526_2192.t3 5.8005
R3831 a_14526_2192.n1 a_14526_2192.t5 5.8005
R3832 a_14526_2192.n0 a_14526_2192.t1 5.8005
R3833 a_14526_2192.n0 a_14526_2192.t0 5.8005
R3834 a_14526_2192.n3 a_14526_2192.t2 5.8005
R3835 a_14526_2192.t4 a_14526_2192.n3 5.8005
R3836 term_6.n1 term_6.t5 734.539
R3837 term_6.n1 term_6.t4 233.26
R3838 term_6.n2 term_6.n1 162.399
R3839 term_6.n2 term_6.n0 75.5108
R3840 term_6.n4 term_6.n3 66.3172
R3841 term_6.n3 term_6.t0 17.4005
R3842 term_6.n3 term_6.t2 17.4005
R3843 term_6.n0 term_6.t3 9.52217
R3844 term_6.n0 term_6.t1 9.52217
R3845 term_6 term_6.n4 5.08746
R3846 term_6.n4 term_6.n2 0.3755
R3847 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 879.481
R3848 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 742.783
R3849 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 665.16
R3850 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 623.388
R3851 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 523.774
R3852 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 431.807
R3853 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 427.875
R3854 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 357.26
R3855 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 208.537
R3856 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 168.077
R3857 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R3858 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R3859 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R3860 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 11.1806
R3861 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R3862 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R3863 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R3864 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R3865 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R3866 term_4.n1 term_4.t5 734.539
R3867 term_4.n1 term_4.t4 233.26
R3868 term_4.n2 term_4.n1 162.399
R3869 term_4.n2 term_4.n0 75.5108
R3870 term_4.n4 term_4.n3 66.3172
R3871 term_4.n3 term_4.t3 17.4005
R3872 term_4.n3 term_4.t0 17.4005
R3873 term_4.n0 term_4.t1 9.52217
R3874 term_4.n0 term_4.t2 9.52217
R3875 term_4 term_4.n4 5.08746
R3876 term_4.n4 term_4.n2 0.3755
R3877 term_2.n1 term_2.t5 734.539
R3878 term_2.n1 term_2.t4 233.26
R3879 term_2.n2 term_2.n1 162.399
R3880 term_2.n2 term_2.n0 75.5108
R3881 term_2.n4 term_2.n3 66.3172
R3882 term_2.n3 term_2.t0 17.4005
R3883 term_2.n3 term_2.t2 17.4005
R3884 term_2.n0 term_2.t3 9.52217
R3885 term_2.n0 term_2.t1 9.52217
R3886 term_2 term_2.n4 5.08746
R3887 term_2.n4 term_2.n2 0.3755
R3888 a_7680_2192.n2 a_7680_2192.n1 34.9195
R3889 a_7680_2192.n2 a_7680_2192.n0 25.5407
R3890 a_7680_2192.n3 a_7680_2192.n2 25.2907
R3891 a_7680_2192.n1 a_7680_2192.t3 5.8005
R3892 a_7680_2192.n1 a_7680_2192.t5 5.8005
R3893 a_7680_2192.n0 a_7680_2192.t1 5.8005
R3894 a_7680_2192.n0 a_7680_2192.t0 5.8005
R3895 a_7680_2192.t4 a_7680_2192.n3 5.8005
R3896 a_7680_2192.n3 a_7680_2192.t2 5.8005
R3897 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 890.727
R3898 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 742.783
R3899 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 665.16
R3900 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 623.388
R3901 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 523.774
R3902 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 431.807
R3903 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 427.875
R3904 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 364.733
R3905 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 208.5
R3906 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 168.007
R3907 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R3908 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 31.2728
R3909 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 31.0337
R3910 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R3911 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R3912 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 9.08234
R3913 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R3914 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R3915 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R3916 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R3917 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R3918 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 879.481
R3919 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 742.783
R3920 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 665.16
R3921 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 623.388
R3922 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 523.774
R3923 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 431.807
R3924 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 427.875
R3925 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 357.26
R3926 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 208.537
R3927 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 168.077
R3928 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R3929 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R3930 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R3931 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 11.1806
R3932 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R3933 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R3934 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R3935 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R3936 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R3937 a_12244_2192.n2 a_12244_2192.n1 34.9195
R3938 a_12244_2192.n2 a_12244_2192.n0 25.5407
R3939 a_12244_2192.n3 a_12244_2192.n2 25.2907
R3940 a_12244_2192.n1 a_12244_2192.t5 5.8005
R3941 a_12244_2192.n1 a_12244_2192.t3 5.8005
R3942 a_12244_2192.n0 a_12244_2192.t1 5.8005
R3943 a_12244_2192.n0 a_12244_2192.t0 5.8005
R3944 a_12244_2192.t4 a_12244_2192.n3 5.8005
R3945 a_12244_2192.n3 a_12244_2192.t2 5.8005
C0 term_5 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.53e-22
C1 stop_strong a_10464_730# 9.87e-20
C2 stop_strong a_12746_730# 9.87e-20
C3 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/delay_unit_2_0.in_2 0.237663f
C4 a_12100_160# a_10502_1376# 0.006618f
C5 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VDD 2.58216f
C6 saff_delay_unit_5/delay_unit_2_0.in_1 VDD 5.0846f
C7 a_12100_160# a_12784_1376# 0.005826f
C8 a_5254_160# saff_delay_unit_2/saff_2_0.nq 0.014786f
C9 a_658_2192# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 1.06381f
C10 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_1 0.868752f
C11 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_2 0.285853f
C12 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.006183f
C13 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_1 0.285853f
C14 saff_delay_unit_1/saff_2_0.nq saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.231514f
C15 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5522_730# 0.003664f
C16 saff_delay_unit_2/saff_2_0.nq VDD 0.712407f
C17 stop_strong a_2940_2192# 4.3e-19
C18 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_5254_160# 3.41e-19
C19 a_3240_296# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.010872f
C20 a_14382_160# a_14650_296# 1.02e-19
C21 a_10086_296# VDD 6.18e-19
C22 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VDD 2.58733f
C23 a_5900_730# saff_delay_unit_2/saff_2_0.nq 0.504416f
C24 a_1374_1376# VDD 1.4126f
C25 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VDD 2.58216f
C26 saff_delay_unit_4/delay_unit_2_0.in_1 a_7804_730# 1.47e-19
C27 a_2972_160# term_1 0.098152f
C28 a_7504_2192# a_7536_160# 2.08e-21
C29 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 term_6 1.53e-22
C30 a_15028_296# VDD 6.18e-19
C31 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C32 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 term_5 0.200954f
C33 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.nq 0.132388f
C34 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.747722f
C35 a_3618_296# VDD 6.18e-19
C36 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/delay_unit_2_0.in_2 0.237663f
C37 a_1336_730# VDD 0.497547f
C38 term_4 VDD 0.589355f
C39 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.99e-19
C40 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_690_160# 0.196687f
C41 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/delay_unit_2_0.in_2 0.018644f
C42 a_1374_1376# a_690_160# 0.005826f
C43 VDD saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 2.44381f
C44 a_9818_160# VDD 1.43296f
C45 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.010157f
C46 saff_delay_unit_2/saff_2_0.nq a_5522_296# 0.005553f
C47 a_14382_160# saff_delay_unit_7/delay_unit_2_0.in_1 3.84e-19
C48 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 9.61e-20
C49 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_2 0.006183f
C50 VDD a_7536_160# 1.43296f
C51 a_3240_730# term_1 0.492009f
C52 saff_delay_unit_1/saff_2_0.nq saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 2.59e-20
C53 a_12100_160# saff_delay_unit_5/saff_2_0.nq 0.014786f
C54 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.nq 0.132388f
C55 a_12100_160# saff_delay_unit_6/delay_unit_2_0.in_1 3.84e-19
C56 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 1.99e-19
C57 saff_delay_unit_6/delay_unit_2_0.in_2 a_12068_2192# 0.007929f
C58 term_3 a_7804_730# 0.492009f
C59 saff_delay_unit_1/saff_2_0.nq a_3618_296# 0.174293f
C60 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.nq 0.132388f
C61 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/delay_unit_2_0.in_2 0.018644f
C62 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.747722f
C63 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/delay_unit_2_0.in_2 0.441403f
C64 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VDD 2.58216f
C65 saff_delay_unit_5/saff_2_0.nq a_12368_730# 0.013457f
C66 a_1374_1376# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 3.22e-19
C67 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 4.28602f
C68 a_17310_296# VDD 6.18e-19
C69 a_12368_730# saff_delay_unit_6/delay_unit_2_0.in_1 1.47e-19
C70 a_7804_296# a_7536_160# 1.02e-19
C71 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_3618_296# 0.012202f
C72 a_2972_160# a_2940_2192# 2.08e-21
C73 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.747722f
C74 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/delay_unit_2_0.in_2 0.237663f
C75 term_3 a_8182_296# 0.005553f
C76 a_958_296# term_0 0.188081f
C77 a_9818_160# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.41e-19
C78 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_2 0.285853f
C79 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.nq 0.231514f
C80 saff_delay_unit_5/saff_2_0.nq a_12368_296# 0.005553f
C81 a_10464_296# a_10502_1376# 1.02e-19
C82 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5254_160# 0.164202f
C83 stop_strong saff_delay_unit_1/delay_unit_2_0.in_1 0.19403f
C84 delay_unit_2_0.out_2 VDD 1.94209f
C85 stop_strong saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.378283f
C86 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C87 a_7536_160# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.196687f
C88 a_15028_296# saff_delay_unit_6/saff_2_0.nq 0.174293f
C89 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/delay_unit_2_0.in_1 0.003768f
C90 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.nq 0.231514f
C91 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.28602f
C92 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5900_730# 0.033952f
C93 a_17310_296# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.012202f
C94 saff_delay_unit_3/delay_unit_2_0.in_2 a_5938_1376# 5.04e-20
C95 saff_delay_unit_5/delay_unit_2_0.in_1 term_4 1.13e-20
C96 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.nq 2.59e-20
C97 stop_strong term_5 7.9e-20
C98 stop_strong term_0 7.9e-20
C99 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/delay_unit_2_0.in_2 0.441403f
C100 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_2 0.961347f
C101 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.138536f
C102 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 3.6e-19
C103 a_9818_160# saff_delay_unit_5/delay_unit_2_0.in_1 3.84e-19
C104 a_1374_1376# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.162437f
C105 start_pos saff_delay_unit_1/delay_unit_2_0.in_1 0.761263f
C106 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_1374_1376# 7.19e-22
C107 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_10502_1376# 3.22e-19
C108 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/delay_unit_2_0.in_1 4.73e-19
C109 a_12784_1376# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.197072f
C110 a_958_296# VDD 6.18e-19
C111 stop_strong a_7504_2192# 4.3e-19
C112 a_10086_296# term_4 0.188081f
C113 a_1336_730# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.003607f
C114 stop_strong saff_delay_unit_2/delay_unit_2_0.in_2 0.538328f
C115 a_1336_730# a_1374_1376# 0.030083f
C116 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_15028_296# 0.012202f
C117 a_10086_296# a_9818_160# 1.02e-19
C118 saff_delay_unit_4/saff_2_0.nq VDD 0.712407f
C119 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 6.79e-20
C120 a_8220_1376# a_8182_296# 1.02e-19
C121 stop_strong a_658_2192# 3.98e-19
C122 saff_delay_unit_2/saff_2_0.nq a_7536_160# 6.08e-20
C123 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.nq 2.59e-20
C124 a_958_296# a_690_160# 1.02e-19
C125 a_15066_1376# VDD 1.4126f
C126 term_6 a_14382_160# 0.098152f
C127 a_7504_2192# saff_delay_unit_4/delay_unit_2_0.in_2 0.007929f
C128 VDD saff_delay_unit_3/saff_2_0.nq 0.712407f
C129 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C130 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C131 term_4 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.105071f
C132 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/delay_unit_2_0.in_1 4.73e-19
C133 start_neg saff_delay_unit_1/delay_unit_2_0.in_1 0.623834f
C134 a_9818_160# term_4 0.098152f
C135 stop_strong VDD 21.0165f
C136 a_9818_160# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.164202f
C137 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.73e-19
C138 term_3 a_8182_730# 0.013457f
C139 a_10464_296# a_10464_730# 0.003413f
C140 stop_strong saff_delay_unit_6/delay_unit_2_0.in_2 0.538328f
C141 stop_strong a_5900_730# 9.87e-20
C142 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_10502_1376# 0.162437f
C143 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12746_296# 0.012202f
C144 a_12784_1376# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.36e-21
C145 a_7804_296# saff_delay_unit_3/saff_2_0.nq 0.005553f
C146 term_2 a_5900_296# 0.005553f
C147 saff_delay_unit_4/delay_unit_2_0.in_2 VDD 3.25148f
C148 a_16932_296# saff_delay_unit_7/saff_2_0.nq 0.005553f
C149 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_15066_1376# 3.22e-19
C150 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.59e-20
C151 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.747722f
C152 term_6 a_14650_296# 0.188081f
C153 saff_delay_unit_5/saff_2_0.nq saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.231514f
C154 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/delay_unit_2_0.in_1 0.138536f
C155 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/saff_2_0.nq 0.231514f
C156 start_pos VDD 2.19021f
C157 a_1336_296# saff_delay_unit_0/saff_2_0.nq 0.174293f
C158 a_12100_160# term_5 0.098152f
C159 stop_strong saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.378271f
C160 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 6.79e-20
C161 saff_delay_unit_3/saff_2_0.nq saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.132388f
C162 stop_strong saff_delay_unit_1/saff_2_0.nq 6.62e-20
C163 term_7 a_17348_1376# 0.014789f
C164 a_17348_1376# a_16664_160# 0.005826f
C165 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.747722f
C166 a_2972_160# saff_delay_unit_2/delay_unit_2_0.in_2 4.55e-19
C167 a_12746_730# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.033952f
C168 stop_strong saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.140412f
C169 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12068_2192# 1.06381f
C170 a_9786_2192# saff_delay_unit_5/delay_unit_2_0.in_1 0.192064f
C171 a_12368_730# term_5 0.492009f
C172 term_6 saff_delay_unit_7/delay_unit_2_0.in_1 1.13e-20
C173 stop_strong saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.378283f
C174 saff_delay_unit_2/delay_unit_2_0.in_1 term_1 1.13e-20
C175 a_8220_1376# a_8182_730# 0.030083f
C176 a_14650_730# a_14382_160# 0.030392f
C177 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_5/delay_unit_2_0.in_1 0.001059f
C178 a_15066_1376# saff_delay_unit_6/saff_2_0.nq 0.100257f
C179 start_neg VDD 1.11527f
C180 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.237663f
C181 term_5 a_12368_296# 0.188081f
C182 a_2972_160# a_3240_296# 1.02e-19
C183 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_8220_1376# 7.19e-22
C184 a_15028_730# VDD 0.497547f
C185 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_15066_1376# 0.162437f
C186 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/delay_unit_2_0.in_2 0.018644f
C187 saff_delay_unit_0/saff_2_0.nq saff_delay_unit_1/delay_unit_2_0.in_1 0.001059f
C188 a_2972_160# VDD 1.43296f
C189 a_958_296# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.010872f
C190 stop_strong saff_delay_unit_6/saff_2_0.nq 6.62e-20
C191 saff_delay_unit_5/saff_2_0.nq saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.59e-20
C192 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_7536_160# 1.15e-21
C193 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/delay_unit_2_0.in_1 0.010157f
C194 stop_strong saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.140412f
C195 a_12100_160# VDD 1.43296f
C196 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_17348_1376# 0.162437f
C197 a_10086_296# saff_delay_unit_4/saff_2_0.nq 0.005553f
C198 stop_strong saff_delay_unit_5/delay_unit_2_0.in_1 0.197172f
C199 VDD saff_delay_unit_7/saff_2_0.nq 0.712407f
C200 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_7804_730# 0.003664f
C201 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_10464_730# 0.003607f
C202 a_12100_160# saff_delay_unit_6/delay_unit_2_0.in_2 4.55e-19
C203 a_9786_2192# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.09966f
C204 a_9786_2192# a_9818_160# 2.08e-21
C205 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_1 0.761263f
C206 stop_strong saff_delay_unit_2/saff_2_0.nq 6.62e-20
C207 saff_delay_unit_0/saff_2_0.nq term_0 0.227882f
C208 a_12784_1376# a_14382_160# 0.006618f
C209 a_3240_296# a_3240_730# 0.003413f
C210 saff_delay_unit_4/saff_2_0.nq term_4 0.227882f
C211 a_14650_730# a_14650_296# 0.003413f
C212 VDD a_10086_730# 0.497771f
C213 a_12368_730# VDD 0.497771f
C214 a_15028_296# a_15066_1376# 1.02e-19
C215 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_1 0.285853f
C216 a_3240_730# VDD 0.497771f
C217 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_2 0.868752f
C218 stop_strong saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.140241f
C219 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_15066_1376# 0.197072f
C220 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.231514f
C221 a_9818_160# saff_delay_unit_4/saff_2_0.nq 0.014786f
C222 stop_strong a_1374_1376# 0.001226f
C223 stop_strong saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.140412f
C224 a_2972_160# saff_delay_unit_1/saff_2_0.nq 0.014786f
C225 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_2 0.019931f
C226 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5222_2192# 1.06381f
C227 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_8182_296# 0.012202f
C228 VDD saff_delay_unit_7/delay_unit_2_0.in_2 3.25148f
C229 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 stop_strong 0.378283f
C230 VDD a_12368_296# 6.18e-19
C231 term_7 a_17310_730# 0.013457f
C232 a_1336_730# stop_strong 9.87e-20
C233 stop_strong term_4 7.9e-20
C234 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_958_730# 0.003664f
C235 a_9818_160# saff_delay_unit_3/saff_2_0.nq 6.08e-20
C236 a_16932_730# saff_delay_unit_7/saff_2_0.nq 0.013457f
C237 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.nq 0.231514f
C238 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_2 0.019931f
C239 saff_delay_unit_2/delay_unit_2_0.in_1 a_2940_2192# 0.192064f
C240 stop_strong saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.378283f
C241 a_2972_160# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.164202f
C242 a_14650_730# saff_delay_unit_7/delay_unit_2_0.in_1 1.47e-19
C243 saff_delay_unit_3/delay_unit_2_0.in_2 a_5254_160# 4.55e-19
C244 a_7536_160# saff_delay_unit_3/saff_2_0.nq 0.014786f
C245 start_pos saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.73e-19
C246 saff_delay_unit_3/delay_unit_2_0.in_2 VDD 3.25148f
C247 stop_strong a_12068_2192# 4.3e-19
C248 saff_delay_unit_1/saff_2_0.nq a_3240_730# 0.013457f
C249 saff_delay_unit_0/saff_2_0.nq VDD 0.712378f
C250 a_15028_730# saff_delay_unit_6/saff_2_0.nq 0.504416f
C251 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_2 0.018644f
C252 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.018644f
C253 saff_delay_unit_5/delay_unit_2_0.in_2 a_10502_1376# 5.04e-20
C254 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_15028_730# 0.003607f
C255 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_15066_1376# 2.36e-21
C256 saff_delay_unit_5/saff_2_0.nq a_14382_160# 6.08e-20
C257 VDD a_7804_730# 0.497771f
C258 a_3240_730# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003664f
C259 saff_delay_unit_4/delay_unit_2_0.in_2 a_7536_160# 4.55e-19
C260 saff_delay_unit_0/saff_2_0.nq a_690_160# 0.014786f
C261 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_17310_730# 0.003607f
C262 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 stop_strong 0.140412f
C263 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.nq 2.59e-20
C264 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 term_5 0.105071f
C265 a_5938_1376# a_5900_296# 1.02e-19
C266 a_2972_160# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 3.41e-19
C267 VDD a_8182_296# 6.18e-19
C268 a_2972_160# a_1374_1376# 0.006618f
C269 a_2972_160# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.196687f
C270 a_7804_296# a_7804_730# 0.003413f
C271 a_10464_296# VDD 6.18e-19
C272 saff_delay_unit_1/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_2 0.961347f
C273 a_15028_296# a_15028_730# 0.003413f
C274 saff_delay_unit_5/delay_unit_2_0.in_1 a_10086_730# 1.47e-19
C275 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_15028_730# 0.033952f
C276 saff_delay_unit_6/saff_2_0.nq saff_delay_unit_7/delay_unit_2_0.in_2 1.23e-19
C277 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.006183f
C278 stop_strong saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.378283f
C279 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_1 4.73e-19
C280 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_8182_730# 0.033952f
C281 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_2 0.237663f
C282 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 9.61e-20
C283 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 6.79e-20
C284 a_7804_730# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.035356f
C285 saff_delay_unit_3/delay_unit_2_0.in_1 a_5222_2192# 0.192064f
C286 a_10086_296# a_10086_730# 0.003413f
C287 saff_delay_unit_1/delay_unit_2_0.in_2 term_0 3.6e-19
C288 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_1 0.761263f
C289 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/delay_unit_2_0.in_2 9.61e-20
C290 a_12100_160# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.15e-21
C291 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_3240_730# 0.035356f
C292 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_2 0.868752f
C293 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C294 term_4 a_10086_730# 0.492009f
C295 a_9786_2192# stop_strong 4.3e-19
C296 a_12100_160# a_12068_2192# 2.08e-21
C297 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_2 0.019931f
C298 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_2 0.441403f
C299 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_1 0.761263f
C300 a_10086_730# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.003664f
C301 a_9818_160# a_10086_730# 0.030392f
C302 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/delay_unit_2_0.in_2 0.441403f
C303 stop_strong saff_delay_unit_4/saff_2_0.nq 6.62e-20
C304 a_658_2192# saff_delay_unit_1/delay_unit_2_0.in_2 0.007929f
C305 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_2/saff_2_0.nq 1.23e-19
C306 term_6 a_14650_730# 0.492009f
C307 stop_strong a_15066_1376# 0.001226f
C308 stop_strong saff_delay_unit_3/saff_2_0.nq 6.62e-20
C309 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12100_160# 0.196687f
C310 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/delay_unit_2_0.in_2 1.17e-19
C311 a_16632_2192# a_16664_160# 2.08e-21
C312 saff_delay_unit_0/saff_2_0.nq saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.132388f
C313 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_2/delay_unit_2_0.in_2 0.961347f
C314 saff_delay_unit_0/saff_2_0.nq a_1374_1376# 0.100257f
C315 saff_delay_unit_1/delay_unit_2_0.in_2 VDD 3.25162f
C316 a_17310_296# saff_delay_unit_7/saff_2_0.nq 0.174293f
C317 VDD a_8182_730# 0.497547f
C318 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 term_2 0.200954f
C319 a_1336_730# saff_delay_unit_0/saff_2_0.nq 0.504416f
C320 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12368_730# 0.035356f
C321 saff_delay_unit_4/delay_unit_2_0.in_2 saff_delay_unit_3/saff_2_0.nq 1.23e-19
C322 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VDD 2.58216f
C323 saff_delay_unit_1/delay_unit_2_0.in_2 a_690_160# 4.55e-19
C324 a_12784_1376# term_6 6.12e-20
C325 stop_strong saff_delay_unit_4/delay_unit_2_0.in_2 0.538328f
C326 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_2 1.17e-19
C327 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/delay_unit_2_0.in_2 1.17e-19
C328 saff_delay_unit_2/delay_unit_2_0.in_1 VDD 5.0846f
C329 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12368_296# 0.010872f
C330 start_pos stop_strong 0.002264f
C331 a_3656_1376# term_2 6.12e-20
C332 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_16632_2192# 1.06381f
C333 a_7804_730# a_7536_160# 0.030392f
C334 a_10464_296# term_4 0.005553f
C335 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 6.79e-20
C336 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/delay_unit_2_0.in_1 7.03e-19
C337 a_14350_2192# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 1.06381f
C338 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/delay_unit_2_0.in_1 0.010157f
C339 a_8182_730# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.003607f
C340 a_17348_1376# VDD 1.41226f
C341 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/delay_unit_2_0.in_2 0.018644f
C342 a_10464_296# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.012202f
C343 a_15066_1376# a_15028_730# 0.030083f
C344 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.6e-19
C345 a_12100_160# saff_delay_unit_4/saff_2_0.nq 6.08e-20
C346 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_1/saff_2_0.nq 0.001059f
C347 start_neg stop_strong 0.005743f
C348 saff_delay_unit_4/delay_unit_2_0.in_1 term_3 1.13e-20
C349 stop_strong a_15028_730# 9.87e-20
C350 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 term_1 1.53e-22
C351 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/delay_unit_2_0.in_2 0.441403f
C352 saff_delay_unit_4/saff_2_0.nq a_10086_730# 0.013457f
C353 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.99e-19
C354 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_14350_2192# 0.09966f
C355 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.138536f
C356 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 term_4 4.1e-22
C357 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/delay_unit_2_0.in_2 9.61e-20
C358 stop_strong saff_delay_unit_7/saff_2_0.nq 6.62e-20
C359 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_17348_1376# 0.197072f
C360 a_5938_1376# term_2 0.014789f
C361 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C362 term_7 a_16664_160# 0.098152f
C363 VDD a_14382_160# 1.43296f
C364 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/delay_unit_2_0.in_1 0.501329f
C365 start_neg start_pos 0.620375f
C366 saff_delay_unit_3/delay_unit_2_0.in_1 term_2 1.13e-20
C367 a_15066_1376# saff_delay_unit_7/delay_unit_2_0.in_2 5.04e-20
C368 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_3656_1376# 7.19e-22
C369 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/delay_unit_2_0.in_2 0.237663f
C370 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_12068_2192# 0.09966f
C371 a_1374_1376# saff_delay_unit_1/delay_unit_2_0.in_2 5.04e-20
C372 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/delay_unit_2_0.in_2 0.006183f
C373 a_958_296# saff_delay_unit_0/saff_2_0.nq 0.005553f
C374 VDD a_5900_296# 6.18e-19
C375 stop_strong saff_delay_unit_7/delay_unit_2_0.in_2 0.538328f
C376 a_10086_296# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.010872f
C377 a_5900_730# a_5900_296# 0.003413f
C378 a_5254_160# a_5222_2192# 2.08e-21
C379 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 4.28602f
C380 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.010157f
C381 VDD a_14650_296# 6.18e-19
C382 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 term_7 0.200954f
C383 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 term_4 0.200954f
C384 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/delay_unit_2_0.in_1 0.501329f
C385 a_17310_730# VDD 0.497547f
C386 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_16664_160# 0.196687f
C387 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_17348_1376# 2.36e-21
C388 a_958_730# saff_delay_unit_1/delay_unit_2_0.in_1 1.47e-19
C389 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 4.28602f
C390 stop_strong saff_delay_unit_3/delay_unit_2_0.in_2 0.538328f
C391 a_9818_160# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.196687f
C392 stop_strong saff_delay_unit_0/saff_2_0.nq 6.62e-20
C393 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_1 0.761263f
C394 a_7804_730# saff_delay_unit_3/saff_2_0.nq 0.013457f
C395 saff_delay_unit_5/delay_unit_2_0.in_2 VDD 3.25148f
C396 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_8220_1376# 2.36e-21
C397 saff_delay_unit_3/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C398 a_10464_296# saff_delay_unit_4/saff_2_0.nq 0.174293f
C399 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5938_1376# 0.162437f
C400 a_958_730# term_0 0.492009f
C401 a_3656_1376# term_1 0.014789f
C402 VDD saff_delay_unit_7/delay_unit_2_0.in_1 5.0846f
C403 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_5/delay_unit_2_0.in_2 0.019931f
C404 a_3618_730# a_3656_1376# 0.030083f
C405 a_14382_160# saff_delay_unit_6/saff_2_0.nq 0.014786f
C406 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_17310_730# 0.033952f
C407 a_12784_1376# a_12746_296# 1.02e-19
C408 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/delay_unit_2_0.in_1 0.501329f
C409 a_8182_296# saff_delay_unit_3/saff_2_0.nq 0.174293f
C410 saff_delay_unit_6/delay_unit_2_0.in_2 saff_delay_unit_7/delay_unit_2_0.in_1 0.868752f
C411 term_3 a_8220_1376# 0.014789f
C412 a_2972_160# a_3240_730# 0.030392f
C413 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.6e-19
C414 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1336_296# 0.012202f
C415 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_14382_160# 0.196687f
C416 a_5938_1376# term_3 6.12e-20
C417 a_12100_160# a_12368_730# 0.030392f
C418 saff_delay_unit_5/saff_2_0.nq a_12784_1376# 0.100257f
C419 a_5522_730# term_2 0.492009f
C420 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_1 7.03e-19
C421 a_12100_160# a_12368_296# 1.02e-19
C422 a_10502_1376# a_10464_730# 0.030083f
C423 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 1.17e-19
C424 a_3618_730# term_1 0.013457f
C425 a_12784_1376# a_12746_730# 0.030083f
C426 saff_delay_unit_6/saff_2_0.nq a_14650_296# 0.005553f
C427 saff_delay_unit_2/saff_2_0.nq a_5900_296# 0.174293f
C428 a_958_730# VDD 0.497771f
C429 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_14382_160# 0.164202f
C430 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/delay_unit_2_0.in_1 7.03e-19
C431 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_14650_296# 0.010872f
C432 a_2972_160# saff_delay_unit_0/saff_2_0.nq 6.08e-20
C433 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 term_2 4.1e-22
C434 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/delay_unit_2_0.in_1 0.138536f
C435 stop_strong saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.378283f
C436 a_17310_296# a_17348_1376# 1.02e-19
C437 a_12368_730# a_12368_296# 0.003413f
C438 a_14350_2192# stop_strong 4.3e-19
C439 a_958_730# a_690_160# 0.030392f
C440 saff_delay_unit_5/saff_2_0.nq a_12746_296# 0.174293f
C441 a_9786_2192# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 1.06381f
C442 saff_delay_unit_6/saff_2_0.nq saff_delay_unit_7/delay_unit_2_0.in_1 0.001059f
C443 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_2 0.961347f
C444 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 term_0 0.105071f
C445 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_1 0.501329f
C446 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.132388f
C447 saff_delay_unit_5/saff_2_0.nq saff_delay_unit_6/delay_unit_2_0.in_1 0.001059f
C448 a_12746_730# a_12746_296# 0.003413f
C449 stop_strong saff_delay_unit_1/delay_unit_2_0.in_2 0.538328f
C450 a_8182_730# saff_delay_unit_3/saff_2_0.nq 0.504416f
C451 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/delay_unit_2_0.in_2 9.61e-20
C452 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/delay_unit_2_0.in_1 0.138536f
C453 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_14382_160# 3.41e-19
C454 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5522_730# 0.035356f
C455 stop_strong a_8182_730# 9.87e-20
C456 saff_delay_unit_5/saff_2_0.nq a_12746_730# 0.504416f
C457 stop_strong saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.140412f
C458 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_658_2192# 0.09966f
C459 term_6 VDD 0.589355f
C460 saff_delay_unit_5/delay_unit_2_0.in_2 term_4 3.6e-19
C461 a_5254_160# term_2 0.098152f
C462 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_1 0.138536f
C463 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.441403f
C464 stop_strong saff_delay_unit_2/delay_unit_2_0.in_1 0.197172f
C465 a_9818_160# saff_delay_unit_5/delay_unit_2_0.in_2 4.55e-19
C466 term_2 VDD 0.589355f
C467 start_pos saff_delay_unit_1/delay_unit_2_0.in_2 0.285853f
C468 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.747722f
C469 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VDD 2.45307f
C470 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/delay_unit_2_0.in_2 0.006183f
C471 a_16932_296# term_7 0.188081f
C472 a_16932_296# a_16664_160# 1.02e-19
C473 a_16632_2192# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.09966f
C474 a_5900_730# term_2 0.013457f
C475 a_7504_2192# saff_delay_unit_4/delay_unit_2_0.in_1 0.192064f
C476 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5900_296# 0.012202f
C477 a_17310_296# a_17310_730# 0.003413f
C478 a_12100_160# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.164202f
C479 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 term_3 0.105071f
C480 term_6 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 4.1e-22
C481 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_690_160# 0.164202f
C482 stop_strong a_17348_1376# 0.001226f
C483 a_958_730# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.035356f
C484 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/delay_unit_2_0.in_2 0.006183f
C485 start_neg saff_delay_unit_1/delay_unit_2_0.in_2 0.019727f
C486 term_2 a_5522_296# 0.188081f
C487 a_12368_730# saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.003664f
C488 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5222_2192# 0.09966f
C489 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.006183f
C490 term_5 a_10502_1376# 6.12e-20
C491 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/delay_unit_2_0.in_1 0.010157f
C492 saff_delay_unit_4/delay_unit_2_0.in_1 VDD 5.0846f
C493 a_12784_1376# term_5 0.014789f
C494 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_2 9.61e-20
C495 a_14350_2192# saff_delay_unit_7/delay_unit_2_0.in_2 0.007929f
C496 a_16932_296# saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.010872f
C497 a_15066_1376# a_14382_160# 0.005826f
C498 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_2 1.53e-22
C499 a_14650_730# VDD 0.497771f
C500 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C501 term_6 saff_delay_unit_6/saff_2_0.nq 0.227882f
C502 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5254_160# 0.196687f
C503 a_12100_160# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.41e-19
C504 saff_delay_unit_2/delay_unit_2_0.in_2 a_3656_1376# 5.04e-20
C505 a_2972_160# saff_delay_unit_2/delay_unit_2_0.in_1 3.84e-19
C506 term_6 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.200954f
C507 saff_delay_unit_3/delay_unit_2_0.in_1 a_5522_730# 1.47e-19
C508 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VDD 2.58216f
C509 term_7 VDD 0.589355f
C510 VDD a_16664_160# 1.43296f
C511 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_8220_1376# 0.197072f
C512 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5900_730# 0.003607f
C513 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_10086_730# 0.035356f
C514 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_5938_1376# 3.22e-19
C515 a_3656_1376# a_5254_160# 0.006618f
C516 term_3 VDD 0.589355f
C517 a_9786_2192# saff_delay_unit_5/delay_unit_2_0.in_2 0.007929f
C518 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.501329f
C519 term_5 a_12746_296# 0.005553f
C520 VDD a_10502_1376# 1.4126f
C521 a_12784_1376# VDD 1.4126f
C522 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/delay_unit_2_0.in_1 7.03e-19
C523 saff_delay_unit_2/saff_2_0.nq term_2 0.227882f
C524 a_3656_1376# VDD 1.4126f
C525 saff_delay_unit_2/delay_unit_2_0.in_1 a_3240_730# 1.47e-19
C526 saff_delay_unit_2/delay_unit_2_0.in_2 term_1 3.6e-19
C527 term_6 a_15028_296# 0.005553f
C528 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 term_6 0.105071f
C529 saff_delay_unit_4/saff_2_0.nq saff_delay_unit_5/delay_unit_2_0.in_2 1.23e-19
C530 a_12784_1376# saff_delay_unit_6/delay_unit_2_0.in_2 5.04e-20
C531 stop_strong a_5222_2192# 4.3e-19
C532 saff_delay_unit_5/saff_2_0.nq term_5 0.227882f
C533 stop_strong a_17310_730# 9.87e-20
C534 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5522_296# 0.010872f
C535 saff_delay_unit_6/delay_unit_2_0.in_1 term_5 1.13e-20
C536 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.28602f
C537 term_7 a_16932_730# 0.492009f
C538 term_7 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.105071f
C539 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1374_1376# 0.197072f
C540 saff_delay_unit_0/saff_2_0.nq saff_delay_unit_1/delay_unit_2_0.in_2 1.23e-19
C541 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 6.79e-20
C542 a_7804_296# term_3 0.188081f
C543 a_16932_730# a_16664_160# 0.030392f
C544 a_17348_1376# saff_delay_unit_7/saff_2_0.nq 0.100257f
C545 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_16664_160# 0.164202f
C546 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.6e-19
C547 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VDD 2.56682f
C548 a_1336_730# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.033952f
C549 stop_strong saff_delay_unit_5/delay_unit_2_0.in_2 0.538328f
C550 a_12746_730# term_5 0.013457f
C551 a_3240_296# term_1 0.188081f
C552 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.79e-20
C553 saff_delay_unit_5/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_1 0.761263f
C554 VDD term_1 0.589355f
C555 stop_strong saff_delay_unit_7/delay_unit_2_0.in_1 0.197172f
C556 a_3618_730# VDD 0.497547f
C557 saff_delay_unit_1/saff_2_0.nq a_3656_1376# 0.100257f
C558 a_14650_730# saff_delay_unit_6/saff_2_0.nq 0.013457f
C559 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_3/delay_unit_2_0.in_2 0.285853f
C560 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_3/delay_unit_2_0.in_1 0.868752f
C561 term_3 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.200954f
C562 a_10502_1376# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.36e-21
C563 a_12746_296# VDD 6.18e-19
C564 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_14650_730# 0.035356f
C565 saff_delay_unit_5/delay_unit_2_0.in_2 saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C566 a_5254_160# a_5938_1376# 0.005826f
C567 a_958_296# a_958_730# 0.003413f
C568 VDD a_8220_1376# 1.4126f
C569 a_3656_1376# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.197072f
C570 saff_delay_unit_6/saff_2_0.nq a_16664_160# 6.08e-20
C571 a_5938_1376# VDD 1.4126f
C572 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 4.28602f
C573 saff_delay_unit_5/saff_2_0.nq VDD 0.712407f
C574 saff_delay_unit_3/delay_unit_2_0.in_1 a_5254_160# 3.84e-19
C575 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_16932_730# 0.035356f
C576 a_8182_730# a_8182_296# 0.003413f
C577 saff_delay_unit_6/delay_unit_2_0.in_1 VDD 5.0846f
C578 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 a_16664_160# 3.41e-19
C579 saff_delay_unit_3/delay_unit_2_0.in_1 VDD 5.0846f
C580 saff_delay_unit_2/delay_unit_2_0.in_2 a_2940_2192# 0.007929f
C581 saff_delay_unit_5/saff_2_0.nq saff_delay_unit_6/delay_unit_2_0.in_2 1.23e-19
C582 a_5900_730# a_5938_1376# 0.030083f
C583 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.nq 0.132388f
C584 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_6/delay_unit_2_0.in_2 0.961347f
C585 saff_delay_unit_1/saff_2_0.nq term_1 0.227882f
C586 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 7.03e-19
C587 a_3618_730# saff_delay_unit_1/saff_2_0.nq 0.504416f
C588 VDD a_10464_730# 0.497547f
C589 a_12746_730# VDD 0.497547f
C590 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_14650_730# 0.003664f
C591 a_12784_1376# saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 7.19e-22
C592 a_14382_160# saff_delay_unit_7/delay_unit_2_0.in_2 4.55e-19
C593 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.6e-19
C594 delay_unit_2_0.out_1 VDD 2.23889f
C595 saff_delay_unit_4/delay_unit_2_0.in_1 a_7536_160# 3.84e-19
C596 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_1 0.105071f
C597 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_2 0.105071f
C598 a_3618_730# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.033952f
C599 a_1336_296# term_0 0.005553f
C600 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 term_7 1.53e-22
C601 a_17310_730# saff_delay_unit_7/saff_2_0.nq 0.504416f
C602 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_16664_160# 1.15e-21
C603 a_8220_1376# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.162437f
C604 a_5938_1376# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 7.19e-22
C605 a_3656_1376# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 2.36e-21
C606 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.747722f
C607 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C608 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_3656_1376# 0.162437f
C609 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 a_12784_1376# 3.22e-19
C610 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.73e-19
C611 a_3656_1376# a_3618_296# 1.02e-19
C612 term_4 a_10502_1376# 0.014789f
C613 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_7536_160# 3.41e-19
C614 term_3 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 4.1e-22
C615 a_10502_1376# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.197072f
C616 a_9818_160# a_10502_1376# 0.005826f
C617 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003768f
C618 saff_delay_unit_1/delay_unit_2_0.in_1 term_0 1.13e-20
C619 term_3 a_7536_160# 0.098152f
C620 term_6 a_15066_1376# 0.014789f
C621 stop_strong a_16632_2192# 4.3e-19
C622 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/delay_unit_2_0.in_1 0.003768f
C623 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 6.79e-20
C624 a_1336_296# VDD 6.18e-19
C625 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 term_1 0.200954f
C626 a_1374_1376# term_1 6.12e-20
C627 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.73e-19
C628 a_17310_296# term_7 0.005553f
C629 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_5/delay_unit_2_0.in_1 0.761263f
C630 a_3618_730# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.003607f
C631 stop_strong term_6 7.9e-20
C632 saff_delay_unit_3/delay_unit_2_0.in_2 a_5222_2192# 0.007929f
C633 saff_delay_unit_7/delay_unit_2_0.in_1 saff_delay_unit_7/delay_unit_2_0.in_2 0.961347f
C634 a_3618_296# term_1 0.005553f
C635 a_5522_730# a_5254_160# 0.030392f
C636 saff_delay_unit_2/delay_unit_2_0.in_1 saff_delay_unit_1/delay_unit_2_0.in_2 0.868752f
C637 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_1/delay_unit_2_0.in_1 0.285853f
C638 a_3618_730# a_3618_296# 0.003413f
C639 a_7504_2192# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.09966f
C640 a_2940_2192# saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.09966f
C641 saff_delay_unit_2/saff_2_0.nq a_5938_1376# 0.100257f
C642 a_5522_730# VDD 0.497771f
C643 stop_strong term_2 7.9e-20
C644 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_10502_1376# 7.19e-22
C645 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12784_1376# 0.162437f
C646 a_658_2192# saff_delay_unit_1/delay_unit_2_0.in_1 0.192064f
C647 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.28602f
C648 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 stop_strong 0.377977f
C649 saff_delay_unit_3/delay_unit_2_0.in_1 saff_delay_unit_2/saff_2_0.nq 0.001059f
C650 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_5938_1376# 2.36e-21
C651 term_4 a_8220_1376# 6.12e-20
C652 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_6/delay_unit_2_0.in_1 7.03e-19
C653 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/delay_unit_2_0.in_1 0.010157f
C654 a_8220_1376# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 3.22e-19
C655 saff_delay_unit_1/delay_unit_2_0.in_1 VDD 5.23339f
C656 a_9818_160# a_8220_1376# 0.006618f
C657 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_3 1.53e-22
C658 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C659 a_16932_296# VDD 6.18e-19
C660 saff_delay_unit_6/delay_unit_2_0.in_1 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.003768f
C661 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_3656_1376# 3.22e-19
C662 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 a_14382_160# 1.15e-21
C663 a_14350_2192# a_14382_160# 2.08e-21
C664 a_8220_1376# a_7536_160# 0.005826f
C665 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_3/saff_2_0.nq 0.001059f
C666 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 start_pos 7.03e-19
C667 term_4 a_10464_730# 0.013457f
C668 a_5522_730# a_5522_296# 0.003413f
C669 saff_delay_unit_1/delay_unit_2_0.in_1 a_690_160# 3.84e-19
C670 a_5938_1376# a_7536_160# 0.006618f
C671 saff_delay_unit_6/delay_unit_2_0.in_1 a_12068_2192# 0.192064f
C672 term_5 VDD 0.589355f
C673 stop_strong saff_delay_unit_4/delay_unit_2_0.in_1 0.197172f
C674 a_10464_730# saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.033952f
C675 VDD term_0 0.589355f
C676 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_2940_2192# 1.06381f
C677 saff_delay_unit_6/delay_unit_2_0.in_2 term_5 3.6e-19
C678 term_6 a_15028_730# 0.013457f
C679 a_16932_296# a_16932_730# 0.003413f
C680 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_3/saff_2_0.nq 2.59e-20
C681 a_690_160# term_0 0.098152f
C682 term_7 a_15066_1376# 6.12e-20
C683 saff_delay_unit_2/delay_unit_2_0.in_2 VDD 3.25148f
C684 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/saff_2_0.nq 0.132388f
C685 saff_delay_unit_4/delay_unit_2_0.in_1 saff_delay_unit_4/delay_unit_2_0.in_2 0.961347f
C686 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_1 4.1e-22
C687 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_6/delay_unit_2_0.in_1 0.501329f
C688 saff_delay_unit_0/saff_2_0.nq a_958_730# 0.013457f
C689 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 start_neg 0.007279f
C690 a_15066_1376# a_16664_160# 0.006618f
C691 saff_delay_unit_4/saff_2_0.nq a_10502_1376# 0.100257f
C692 stop_strong saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.140412f
C693 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.28602f
C694 stop_strong term_7 7.9e-20
C695 a_2972_160# saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 1.15e-21
C696 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_1/delay_unit_2_0.in_1 7.03e-19
C697 term_3 saff_delay_unit_3/saff_2_0.nq 0.227882f
C698 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 a_12746_730# 0.003607f
C699 a_5254_160# VDD 1.43296f
C700 a_3240_296# VDD 6.18e-19
C701 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5938_1376# 0.197072f
C702 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/delay_unit_2_0.in_2 0.018644f
C703 stop_strong term_3 7.9e-20
C704 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_4/delay_unit_2_0.in_2 1.17e-19
C705 a_1336_296# a_1374_1376# 1.02e-19
C706 stop_strong a_10502_1376# 0.001226f
C707 a_658_2192# a_690_160# 2.08e-21
C708 stop_strong a_12784_1376# 0.001226f
C709 a_5522_730# saff_delay_unit_2/saff_2_0.nq 0.013457f
C710 stop_strong a_3656_1376# 0.001226f
C711 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_3/delay_unit_2_0.in_1 0.138536f
C712 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_7/delay_unit_2_0.in_1 0.003768f
C713 a_14350_2192# saff_delay_unit_7/delay_unit_2_0.in_1 0.192064f
C714 term_6 saff_delay_unit_7/delay_unit_2_0.in_2 3.6e-19
C715 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_0 4.1e-22
C716 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_1/saff_2_0.nq 1.23e-19
C717 a_1336_730# a_1336_296# 0.003413f
C718 saff_delay_unit_6/delay_unit_2_0.in_2 VDD 3.25148f
C719 a_5900_730# VDD 0.497547f
C720 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_5/delay_unit_2_0.in_1 0.003768f
C721 saff_delay_unit_4/delay_unit_2_0.in_2 term_3 3.6e-19
C722 a_7504_2192# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 1.06381f
C723 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_15066_1376# 7.19e-22
C724 VDD a_690_160# 1.43261f
C725 delay_unit_2_0.out_2 delay_unit_2_0.out_1 0.031607f
C726 a_7804_296# VDD 6.18e-19
C727 stop_strong saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.140399f
C728 a_5254_160# a_5522_296# 1.02e-19
C729 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.441403f
C730 saff_delay_unit_1/saff_2_0.nq a_5254_160# 6.08e-20
C731 a_3240_296# saff_delay_unit_1/saff_2_0.nq 0.005553f
C732 a_16932_730# VDD 0.497771f
C733 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/delay_unit_2_0.in_1 0.501329f
C734 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C735 VDD a_5522_296# 6.18e-19
C736 saff_delay_unit_1/saff_2_0.nq VDD 0.712407f
C737 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_1/delay_unit_2_0.in_1 4.73e-19
C738 stop_strong term_1 7.9e-20
C739 a_3618_730# stop_strong 9.87e-20
C740 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 saff_delay_unit_5/delay_unit_2_0.in_2 0.237663f
C741 saff_delay_unit_3/delay_unit_2_0.in_2 term_2 3.6e-19
C742 a_8220_1376# saff_delay_unit_3/saff_2_0.nq 0.100257f
C743 VDD saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.58216f
C744 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_5254_160# 1.15e-21
C745 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 term_4 1.53e-22
C746 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_0/saff_2_0.nq 0.231514f
C747 stop_strong a_8220_1376# 0.001226f
C748 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 term_0 0.200954f
C749 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VDD 2.44381f
C750 saff_delay_unit_4/saff_2_0.nq a_10464_730# 0.504416f
C751 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C752 a_9818_160# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.15e-21
C753 a_1374_1376# term_0 0.014789f
C754 saff_delay_unit_5/saff_2_0.nq stop_strong 6.62e-20
C755 stop_strong a_5938_1376# 0.001226f
C756 stop_strong saff_delay_unit_6/delay_unit_2_0.in_1 0.197172f
C757 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 term_5 4.1e-22
C758 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_16932_730# 0.003664f
C759 a_17348_1376# a_17310_730# 0.030083f
C760 stop_strong saff_delay_unit_3/delay_unit_2_0.in_1 0.197172f
C761 a_1336_730# term_0 0.013457f
C762 term_7 saff_delay_unit_7/saff_2_0.nq 0.227882f
C763 a_7804_296# saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.010872f
C764 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_7536_160# 0.164202f
C765 a_16664_160# saff_delay_unit_7/saff_2_0.nq 0.014786f
C766 VDD saff_delay_unit_6/saff_2_0.nq 0.712407f
C767 a_2972_160# a_3656_1376# 0.005826f
C768 saff_delay_unit_2/delay_unit_2_0.in_2 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 1.17e-19
C769 saff_delay_unit_4/delay_unit_2_0.in_2 a_8220_1376# 5.04e-20
C770 term_7 VSS 0.725415f
C771 term_6 VSS 0.725414f
C772 term_5 VSS 0.725414f
C773 term_4 VSS 0.725414f
C774 term_3 VSS 0.725414f
C775 term_2 VSS 0.725414f
C776 term_1 VSS 0.725414f
C777 term_0 VSS 0.725444f
C778 stop_strong VSS 21.447275f
C779 start_pos VSS 1.197805f
C780 start_neg VSS 1.52205f
C781 VDD VSS 0.140384p
C782 a_17310_296# VSS 0.192064f
C783 a_16932_296# VSS 0.190559f
C784 a_15028_296# VSS 0.192064f
C785 a_17310_730# VSS 0.023462f
C786 a_16932_730# VSS 0.024712f
C787 a_17348_1376# VSS 0.825208f
C788 saff_delay_unit_7/saff_2_0.nq VSS 0.591638f
C789 a_16664_160# VSS 0.82289f
C790 a_14650_296# VSS 0.190559f
C791 a_12746_296# VSS 0.192064f
C792 a_15028_730# VSS 0.023462f
C793 a_14650_730# VSS 0.024712f
C794 a_15066_1376# VSS 0.817309f
C795 saff_delay_unit_6/saff_2_0.nq VSS 0.591435f
C796 a_14382_160# VSS 0.82289f
C797 a_12368_296# VSS 0.190559f
C798 a_10464_296# VSS 0.192064f
C799 a_12746_730# VSS 0.023462f
C800 a_12368_730# VSS 0.024712f
C801 a_12784_1376# VSS 0.817309f
C802 saff_delay_unit_5/saff_2_0.nq VSS 0.591435f
C803 a_12100_160# VSS 0.82289f
C804 a_10086_296# VSS 0.190559f
C805 a_8182_296# VSS 0.192064f
C806 a_10464_730# VSS 0.023462f
C807 a_10086_730# VSS 0.024712f
C808 a_10502_1376# VSS 0.817309f
C809 saff_delay_unit_4/saff_2_0.nq VSS 0.591435f
C810 a_9818_160# VSS 0.82289f
C811 a_7804_296# VSS 0.190559f
C812 a_5900_296# VSS 0.192064f
C813 a_8182_730# VSS 0.023462f
C814 a_7804_730# VSS 0.024712f
C815 a_8220_1376# VSS 0.817309f
C816 saff_delay_unit_3/saff_2_0.nq VSS 0.591435f
C817 a_7536_160# VSS 0.82289f
C818 a_5522_296# VSS 0.190559f
C819 a_3618_296# VSS 0.192064f
C820 a_5900_730# VSS 0.023462f
C821 a_5522_730# VSS 0.024712f
C822 a_5938_1376# VSS 0.817309f
C823 saff_delay_unit_2/saff_2_0.nq VSS 0.591435f
C824 a_5254_160# VSS 0.82289f
C825 a_3240_296# VSS 0.190559f
C826 a_1336_296# VSS 0.192204f
C827 a_3618_730# VSS 0.023462f
C828 a_3240_730# VSS 0.024712f
C829 a_3656_1376# VSS 0.817309f
C830 saff_delay_unit_1/saff_2_0.nq VSS 0.591435f
C831 a_2972_160# VSS 0.82289f
C832 a_958_296# VSS 0.190808f
C833 a_1336_730# VSS 0.023462f
C834 a_958_730# VSS 0.024712f
C835 a_1374_1376# VSS 0.817492f
C836 saff_delay_unit_0/saff_2_0.nq VSS 0.591989f
C837 a_690_160# VSS 0.832702f
C838 a_16632_2192# VSS 0.354057f
C839 a_14350_2192# VSS 0.354057f
C840 a_12068_2192# VSS 0.354057f
C841 a_9786_2192# VSS 0.354057f
C842 a_7504_2192# VSS 0.354057f
C843 a_5222_2192# VSS 0.354057f
C844 a_2940_2192# VSS 0.354057f
C845 a_658_2192# VSS 0.354057f
C846 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VSS 6.497441f
C847 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VSS 6.455006f
C848 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C849 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C850 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C851 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C852 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C853 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C854 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C855 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C856 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C857 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C858 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VSS 6.036491f
C859 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VSS 6.455515f
C860 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VSS 6.037781f
C861 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VSS 7.144324f
C862 delay_unit_2_0.out_2 VSS 1.24762f
C863 delay_unit_2_0.out_1 VSS 0.976728f
C864 saff_delay_unit_7/delay_unit_2_0.in_2 VSS 6.101376f
C865 saff_delay_unit_7/delay_unit_2_0.in_1 VSS 5.6853f
C866 saff_delay_unit_6/delay_unit_2_0.in_2 VSS 6.049282f
C867 saff_delay_unit_6/delay_unit_2_0.in_1 VSS 5.495615f
C868 saff_delay_unit_5/delay_unit_2_0.in_2 VSS 6.049282f
C869 saff_delay_unit_5/delay_unit_2_0.in_1 VSS 5.495615f
C870 saff_delay_unit_4/delay_unit_2_0.in_2 VSS 6.101376f
C871 saff_delay_unit_4/delay_unit_2_0.in_1 VSS 5.495615f
C872 saff_delay_unit_3/delay_unit_2_0.in_2 VSS 6.049282f
C873 saff_delay_unit_3/delay_unit_2_0.in_1 VSS 5.6853f
C874 saff_delay_unit_2/delay_unit_2_0.in_2 VSS 6.101376f
C875 saff_delay_unit_2/delay_unit_2_0.in_1 VSS 5.6853f
C876 saff_delay_unit_1/delay_unit_2_0.in_2 VSS 6.049312f
C877 saff_delay_unit_1/delay_unit_2_0.in_1 VSS 5.644661f
C878 a_12244_2192.t2 VSS 0.059028f
C879 a_12244_2192.t1 VSS 0.059028f
C880 a_12244_2192.t0 VSS 0.059028f
C881 a_12244_2192.n0 VSS 0.139449f
C882 a_12244_2192.t5 VSS 0.059028f
C883 a_12244_2192.t3 VSS 0.059028f
C884 a_12244_2192.n1 VSS 0.258102f
C885 a_12244_2192.n2 VSS 1.11221f
C886 a_12244_2192.n3 VSS 0.136068f
C887 a_12244_2192.t4 VSS 0.059028f
C888 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C889 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C890 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.087567f
C891 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.039891f
C892 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C893 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C894 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.054262f
C895 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.115133f
C896 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C897 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.095888f
C898 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.041221f
C899 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.116123f
C900 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.108538f
C901 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.081767f
C902 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.090596f
C903 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.106694f
C904 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C905 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C906 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.096169f
C907 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.041341f
C908 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C909 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C910 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C911 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C912 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.202807f
C913 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.200111f
C914 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.087824f
C915 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.040008f
C916 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C917 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C918 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C919 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C920 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.107599f
C921 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C922 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.082007f
C923 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.090862f
C924 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C925 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C926 a_7680_2192.t2 VSS 0.059028f
C927 a_7680_2192.t1 VSS 0.059028f
C928 a_7680_2192.t0 VSS 0.059028f
C929 a_7680_2192.n0 VSS 0.139449f
C930 a_7680_2192.t3 VSS 0.059028f
C931 a_7680_2192.t5 VSS 0.059028f
C932 a_7680_2192.n1 VSS 0.258102f
C933 a_7680_2192.n2 VSS 1.11221f
C934 a_7680_2192.n3 VSS 0.136068f
C935 a_7680_2192.t4 VSS 0.059028f
C936 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.774729f
C937 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.95016f
C938 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.088874f
C939 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.040486f
C940 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.099002f
C941 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.204745f
C942 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.055072f
C943 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.055072f
C944 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116852f
C945 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.097319f
C946 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.041836f
C947 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.117856f
C948 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.110158f
C949 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.082987f
C950 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.091949f
C951 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.108286f
C952 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.204745f
C953 saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.765006f
C954 a_14526_2192.t2 VSS 0.059028f
C955 a_14526_2192.t1 VSS 0.059028f
C956 a_14526_2192.t0 VSS 0.059028f
C957 a_14526_2192.n0 VSS 0.139449f
C958 a_14526_2192.t3 VSS 0.059028f
C959 a_14526_2192.t5 VSS 0.059028f
C960 a_14526_2192.n1 VSS 0.258102f
C961 a_14526_2192.n2 VSS 1.11221f
C962 a_14526_2192.n3 VSS 0.136068f
C963 a_14526_2192.t4 VSS 0.059028f
C964 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.096169f
C965 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.041341f
C966 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C967 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C968 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C969 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C970 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.202807f
C971 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C972 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.087824f
C973 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.040008f
C974 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C975 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C976 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C977 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C978 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.107599f
C979 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C980 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.082007f
C981 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.090862f
C982 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C983 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C984 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C985 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.087824f
C986 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.040008f
C987 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C988 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C989 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.202807f
C990 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.096169f
C991 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.041341f
C992 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C993 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.082007f
C994 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.090862f
C995 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C996 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C997 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.107599f
C998 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C999 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C1000 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C1001 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C1002 saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
C1003 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.936187f
C1004 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.087567f
C1005 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.039891f
C1006 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.097546f
C1007 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C1008 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C1009 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.115133f
C1010 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1011 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.095888f
C1012 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.041221f
C1013 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C1014 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.108538f
C1015 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.081767f
C1016 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.090596f
C1017 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C1018 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.398296f
C1019 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.36504f
C1020 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C1021 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 VSS 0.753756f
C1022 a_9698_2192.t6 VSS 0.024913f
C1023 a_9698_2192.t4 VSS 0.024913f
C1024 a_9698_2192.t7 VSS 0.024913f
C1025 a_9698_2192.n0 VSS 0.060272f
C1026 a_9698_2192.t9 VSS 0.024913f
C1027 a_9698_2192.t3 VSS 0.024913f
C1028 a_9698_2192.n1 VSS 0.060114f
C1029 a_9698_2192.t1 VSS 0.024913f
C1030 a_9698_2192.t12 VSS 0.024913f
C1031 a_9698_2192.n2 VSS 0.060114f
C1032 a_9698_2192.t10 VSS 0.024913f
C1033 a_9698_2192.t0 VSS 0.024913f
C1034 a_9698_2192.n3 VSS 0.060114f
C1035 a_9698_2192.t2 VSS 0.097139f
C1036 a_9698_2192.n4 VSS 0.369186f
C1037 a_9698_2192.n5 VSS 0.182473f
C1038 a_9698_2192.n6 VSS 0.22019f
C1039 a_9698_2192.t5 VSS 0.024913f
C1040 a_9698_2192.t11 VSS 0.024913f
C1041 a_9698_2192.n7 VSS 0.052659f
C1042 a_9698_2192.n8 VSS 0.140942f
C1043 a_9698_2192.n9 VSS 0.340434f
C1044 a_9698_2192.n10 VSS 0.057409f
C1045 a_9698_2192.t8 VSS 0.024913f
C1046 a_9962_2192.t5 VSS 0.059028f
C1047 a_9962_2192.t2 VSS 0.059028f
C1048 a_9962_2192.t3 VSS 0.059028f
C1049 a_9962_2192.n0 VSS 0.136068f
C1050 a_9962_2192.t0 VSS 0.059028f
C1051 a_9962_2192.t1 VSS 0.059028f
C1052 a_9962_2192.n1 VSS 0.258102f
C1053 a_9962_2192.n2 VSS 1.11221f
C1054 a_9962_2192.n3 VSS 0.139449f
C1055 a_9962_2192.t4 VSS 0.059028f
C1056 saff_delay_unit_6/delay_unit_2_0.in_1.t10 VSS 0.059113f
C1057 saff_delay_unit_6/delay_unit_2_0.in_1.t13 VSS 0.018532f
C1058 saff_delay_unit_6/delay_unit_2_0.in_1.n0 VSS 0.043408f
C1059 saff_delay_unit_6/delay_unit_2_0.in_1.t18 VSS 0.059113f
C1060 saff_delay_unit_6/delay_unit_2_0.in_1.t8 VSS 0.018532f
C1061 saff_delay_unit_6/delay_unit_2_0.in_1.n1 VSS 0.04376f
C1062 saff_delay_unit_6/delay_unit_2_0.in_1.n2 VSS 0.01701f
C1063 saff_delay_unit_6/delay_unit_2_0.in_1.t12 VSS 0.059113f
C1064 saff_delay_unit_6/delay_unit_2_0.in_1.t15 VSS 0.018532f
C1065 saff_delay_unit_6/delay_unit_2_0.in_1.n3 VSS 0.04376f
C1066 saff_delay_unit_6/delay_unit_2_0.in_1.t17 VSS 0.059113f
C1067 saff_delay_unit_6/delay_unit_2_0.in_1.t19 VSS 0.018532f
C1068 saff_delay_unit_6/delay_unit_2_0.in_1.n4 VSS 0.043408f
C1069 saff_delay_unit_6/delay_unit_2_0.in_1.n5 VSS 0.016864f
C1070 saff_delay_unit_6/delay_unit_2_0.in_1.n6 VSS 0.348947f
C1071 saff_delay_unit_6/delay_unit_2_0.in_1.t0 VSS 0.04785f
C1072 saff_delay_unit_6/delay_unit_2_0.in_1.t1 VSS 0.144836f
C1073 saff_delay_unit_6/delay_unit_2_0.in_1.n7 VSS 0.367599f
C1074 saff_delay_unit_6/delay_unit_2_0.in_1.n8 VSS 0.189684f
C1075 saff_delay_unit_6/delay_unit_2_0.in_1.t3 VSS 0.013076f
C1076 saff_delay_unit_6/delay_unit_2_0.in_1.t2 VSS 0.013076f
C1077 saff_delay_unit_6/delay_unit_2_0.in_1.n9 VSS 0.030628f
C1078 saff_delay_unit_6/delay_unit_2_0.in_1.t7 VSS 0.039228f
C1079 saff_delay_unit_6/delay_unit_2_0.in_1.t6 VSS 0.039228f
C1080 saff_delay_unit_6/delay_unit_2_0.in_1.n10 VSS 0.079915f
C1081 saff_delay_unit_6/delay_unit_2_0.in_1.n11 VSS 0.332497f
C1082 saff_delay_unit_6/delay_unit_2_0.in_1.t14 VSS 0.061404f
C1083 saff_delay_unit_6/delay_unit_2_0.in_1.t9 VSS 0.061404f
C1084 saff_delay_unit_6/delay_unit_2_0.in_1.n12 VSS 0.069322f
C1085 saff_delay_unit_6/delay_unit_2_0.in_1.t11 VSS 0.061404f
C1086 saff_delay_unit_6/delay_unit_2_0.in_1.t16 VSS 0.061404f
C1087 saff_delay_unit_6/delay_unit_2_0.in_1.n13 VSS 0.068946f
C1088 saff_delay_unit_6/delay_unit_2_0.in_1.n14 VSS 0.629493f
C1089 saff_delay_unit_6/delay_unit_2_0.in_1.t4 VSS 0.045922f
C1090 saff_delay_unit_6/delay_unit_2_0.in_1.n15 VSS 0.158606f
C1091 saff_delay_unit_6/delay_unit_2_0.in_1.t5 VSS 0.144836f
C1092 saff_delay_unit_6/delay_unit_2_0.in_1.n16 VSS 0.240372f
C1093 saff_delay_unit_6/delay_unit_2_0.in_1.n17 VSS 0.180663f
C1094 delay_unit_2_0.out_1.t0 VSS 0.020532f
C1095 delay_unit_2_0.out_1.t1 VSS 0.020532f
C1096 delay_unit_2_0.out_1.n0 VSS 0.048092f
C1097 delay_unit_2_0.out_1.t4 VSS 0.061597f
C1098 delay_unit_2_0.out_1.t5 VSS 0.061597f
C1099 delay_unit_2_0.out_1.n1 VSS 0.125485f
C1100 delay_unit_2_0.out_1.n2 VSS 0.522094f
C1101 delay_unit_2_0.out_1.t2 VSS 0.075157f
C1102 delay_unit_2_0.out_1.t3 VSS 0.227425f
C1103 delay_unit_2_0.out_1.n3 VSS 0.55466f
C1104 delay_unit_2_0.out_1.n4 VSS 0.283681f
C1105 delay_unit_2_0.in_2 VSS 0.191069f
C1106 saff_delay_unit_7/saff_2_0.nd.t17 VSS 0.04604f
C1107 saff_delay_unit_7/saff_2_0.nd.t12 VSS 0.04604f
C1108 saff_delay_unit_7/saff_2_0.nd.n0 VSS 0.053939f
C1109 saff_delay_unit_7/saff_2_0.nd.t10 VSS 0.04604f
C1110 saff_delay_unit_7/saff_2_0.nd.t18 VSS 0.04604f
C1111 saff_delay_unit_7/saff_2_0.nd.n1 VSS 0.053696f
C1112 saff_delay_unit_7/saff_2_0.nd.n2 VSS 0.492134f
C1113 saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd VSS 0.376377f
C1114 saff_delay_unit_7/saff_2_0.nd.t19 VSS 0.03874f
C1115 saff_delay_unit_7/saff_2_0.nd.t9 VSS 0.012145f
C1116 saff_delay_unit_7/saff_2_0.nd.n3 VSS 0.028678f
C1117 saff_delay_unit_7/saff_2_0.nd.t14 VSS 0.03874f
C1118 saff_delay_unit_7/saff_2_0.nd.t16 VSS 0.012145f
C1119 saff_delay_unit_7/saff_2_0.nd.n4 VSS 0.028448f
C1120 saff_delay_unit_7/saff_2_0.nd.n5 VSS 0.011146f
C1121 saff_delay_unit_7/saff_2_0.nd.t8 VSS 0.03874f
C1122 saff_delay_unit_7/saff_2_0.nd.t13 VSS 0.012145f
C1123 saff_delay_unit_7/saff_2_0.nd.n6 VSS 0.028678f
C1124 saff_delay_unit_7/saff_2_0.nd.t11 VSS 0.03874f
C1125 saff_delay_unit_7/saff_2_0.nd.t15 VSS 0.012145f
C1126 saff_delay_unit_7/saff_2_0.nd.n7 VSS 0.028448f
C1127 saff_delay_unit_7/saff_2_0.nd.n8 VSS 0.011052f
C1128 saff_delay_unit_7/saff_2_0.nd.n9 VSS 0.134546f
C1129 saff_delay_unit_7/saff_2_0.nd.t7 VSS 0.097382f
C1130 saff_delay_unit_7/saff_2_0.nd.t6 VSS 0.030095f
C1131 saff_delay_unit_7/saff_2_0.nd.n10 VSS 0.266165f
C1132 saff_delay_unit_7/saff_2_0.nd.n11 VSS 0.122739f
C1133 saff_delay_unit_7/saff_2_0.nd.t3 VSS 0.025709f
C1134 saff_delay_unit_7/saff_2_0.nd.t5 VSS 0.025709f
C1135 saff_delay_unit_7/saff_2_0.nd.n12 VSS 0.054977f
C1136 saff_delay_unit_7/saff_2_0.nd.t1 VSS 0.008569f
C1137 saff_delay_unit_7/saff_2_0.nd.t0 VSS 0.008569f
C1138 saff_delay_unit_7/saff_2_0.nd.n13 VSS 0.018604f
C1139 saff_delay_unit_7/saff_2_0.nd.n14 VSS 0.221085f
C1140 saff_delay_unit_7/saff_2_0.nd.t4 VSS 0.097382f
C1141 saff_delay_unit_7/saff_2_0.nd.t2 VSS 0.030095f
C1142 saff_delay_unit_7/saff_2_0.nd.n15 VSS 0.234034f
C1143 saff_delay_unit_7/saff_2_0.nd.n16 VSS 0.050515f
C1144 saff_delay_unit_7/delay_unit_2_0.out_2 VSS 0.082456f
C1145 a_7416_2192.t5 VSS 0.024913f
C1146 a_7416_2192.t4 VSS 0.024913f
C1147 a_7416_2192.t7 VSS 0.024913f
C1148 a_7416_2192.n0 VSS 0.060272f
C1149 a_7416_2192.t10 VSS 0.024913f
C1150 a_7416_2192.t0 VSS 0.024913f
C1151 a_7416_2192.n1 VSS 0.060114f
C1152 a_7416_2192.t2 VSS 0.024913f
C1153 a_7416_2192.t11 VSS 0.024913f
C1154 a_7416_2192.n2 VSS 0.060114f
C1155 a_7416_2192.t12 VSS 0.024913f
C1156 a_7416_2192.t1 VSS 0.024913f
C1157 a_7416_2192.n3 VSS 0.060114f
C1158 a_7416_2192.t3 VSS 0.097139f
C1159 a_7416_2192.n4 VSS 0.369186f
C1160 a_7416_2192.n5 VSS 0.182473f
C1161 a_7416_2192.n6 VSS 0.22019f
C1162 a_7416_2192.t6 VSS 0.024913f
C1163 a_7416_2192.t9 VSS 0.024913f
C1164 a_7416_2192.n7 VSS 0.052659f
C1165 a_7416_2192.n8 VSS 0.140942f
C1166 a_7416_2192.n9 VSS 0.340434f
C1167 a_7416_2192.n10 VSS 0.057409f
C1168 a_7416_2192.t8 VSS 0.024913f
C1169 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C1170 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.096169f
C1171 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.041341f
C1172 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.116331f
C1173 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1174 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C1175 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.114315f
C1176 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.202807f
C1177 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C1178 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.087824f
C1179 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.040008f
C1180 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.097717f
C1181 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.382243f
C1182 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.107599f
C1183 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C1184 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.082007f
C1185 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.090862f
C1186 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.108213f
C1187 saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 VSS 1.24645f
C1188 saff_delay_unit_6/delay_unit_2_0.in_2.t12 VSS 0.039951f
C1189 saff_delay_unit_6/delay_unit_2_0.in_2.t16 VSS 0.012525f
C1190 saff_delay_unit_6/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1191 saff_delay_unit_6/delay_unit_2_0.in_2.t18 VSS 0.039951f
C1192 saff_delay_unit_6/delay_unit_2_0.in_2.t8 VSS 0.012525f
C1193 saff_delay_unit_6/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1194 saff_delay_unit_6/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1195 saff_delay_unit_6/delay_unit_2_0.in_2.t9 VSS 0.039951f
C1196 saff_delay_unit_6/delay_unit_2_0.in_2.t13 VSS 0.012525f
C1197 saff_delay_unit_6/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1198 saff_delay_unit_6/delay_unit_2_0.in_2.t11 VSS 0.039951f
C1199 saff_delay_unit_6/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1200 saff_delay_unit_6/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1201 saff_delay_unit_6/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1202 saff_delay_unit_6/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1203 saff_delay_unit_6/delay_unit_2_0.in_2.t7 VSS 0.100425f
C1204 saff_delay_unit_6/delay_unit_2_0.in_2.t0 VSS 0.031036f
C1205 saff_delay_unit_6/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1206 saff_delay_unit_6/delay_unit_2_0.in_2.t10 VSS 0.047479f
C1207 saff_delay_unit_6/delay_unit_2_0.in_2.t17 VSS 0.047479f
C1208 saff_delay_unit_6/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1209 saff_delay_unit_6/delay_unit_2_0.in_2.t14 VSS 0.047479f
C1210 saff_delay_unit_6/delay_unit_2_0.in_2.t19 VSS 0.047479f
C1211 saff_delay_unit_6/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1212 saff_delay_unit_6/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1213 saff_delay_unit_6/delay_unit_2_0.in_2.t6 VSS 0.026512f
C1214 saff_delay_unit_6/delay_unit_2_0.in_2.t5 VSS 0.026512f
C1215 saff_delay_unit_6/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1216 saff_delay_unit_6/delay_unit_2_0.in_2.t1 VSS 0.008837f
C1217 saff_delay_unit_6/delay_unit_2_0.in_2.t3 VSS 0.008837f
C1218 saff_delay_unit_6/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1219 saff_delay_unit_6/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1220 saff_delay_unit_6/delay_unit_2_0.in_2.t4 VSS 0.100425f
C1221 saff_delay_unit_6/delay_unit_2_0.in_2.t2 VSS 0.031036f
C1222 saff_delay_unit_6/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1223 saff_delay_unit_6/delay_unit_2_0.in_2.n15 VSS 0.052094f
C1224 saff_delay_unit_6/delay_unit_2_0.in_2.n16 VSS 0.126574f
C1225 saff_delay_unit_7/delay_unit_2_0.in_2.t19 VSS 0.039951f
C1226 saff_delay_unit_7/delay_unit_2_0.in_2.t8 VSS 0.012525f
C1227 saff_delay_unit_7/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1228 saff_delay_unit_7/delay_unit_2_0.in_2.t12 VSS 0.039951f
C1229 saff_delay_unit_7/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1230 saff_delay_unit_7/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1231 saff_delay_unit_7/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1232 saff_delay_unit_7/delay_unit_2_0.in_2.t14 VSS 0.039951f
C1233 saff_delay_unit_7/delay_unit_2_0.in_2.t16 VSS 0.012525f
C1234 saff_delay_unit_7/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1235 saff_delay_unit_7/delay_unit_2_0.in_2.t9 VSS 0.039951f
C1236 saff_delay_unit_7/delay_unit_2_0.in_2.t13 VSS 0.012525f
C1237 saff_delay_unit_7/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1238 saff_delay_unit_7/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1239 saff_delay_unit_7/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1240 saff_delay_unit_7/delay_unit_2_0.in_2.t2 VSS 0.100425f
C1241 saff_delay_unit_7/delay_unit_2_0.in_2.t1 VSS 0.031036f
C1242 saff_delay_unit_7/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1243 saff_delay_unit_7/delay_unit_2_0.in_2.t17 VSS 0.047479f
C1244 saff_delay_unit_7/delay_unit_2_0.in_2.t10 VSS 0.047479f
C1245 saff_delay_unit_7/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1246 saff_delay_unit_7/delay_unit_2_0.in_2.t18 VSS 0.047479f
C1247 saff_delay_unit_7/delay_unit_2_0.in_2.t11 VSS 0.047479f
C1248 saff_delay_unit_7/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1249 saff_delay_unit_7/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1250 saff_delay_unit_7/delay_unit_2_0.in_2.t4 VSS 0.026512f
C1251 saff_delay_unit_7/delay_unit_2_0.in_2.t6 VSS 0.026512f
C1252 saff_delay_unit_7/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1253 saff_delay_unit_7/delay_unit_2_0.in_2.t7 VSS 0.008837f
C1254 saff_delay_unit_7/delay_unit_2_0.in_2.t3 VSS 0.008837f
C1255 saff_delay_unit_7/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1256 saff_delay_unit_7/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1257 saff_delay_unit_7/delay_unit_2_0.in_2.t5 VSS 0.100425f
C1258 saff_delay_unit_7/delay_unit_2_0.in_2.t0 VSS 0.031036f
C1259 saff_delay_unit_7/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1260 saff_delay_unit_7/delay_unit_2_0.in_2.n15 VSS 0.126574f
C1261 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.096169f
C1262 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.041341f
C1263 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C1264 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1265 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C1266 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C1267 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.202807f
C1268 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.087824f
C1269 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.040008f
C1270 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C1271 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.200111f
C1272 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C1273 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C1274 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C1275 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.107599f
C1276 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C1277 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.082007f
C1278 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.090862f
C1279 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C1280 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C1281 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1282 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1283 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.087567f
C1284 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.039891f
C1285 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1286 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.201734f
C1287 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1288 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.095888f
C1289 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.041221f
C1290 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C1291 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.108538f
C1292 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.081767f
C1293 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.090596f
C1294 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C1295 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C1296 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C1297 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C1298 saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1299 a_5398_2192.t2 VSS 0.059028f
C1300 a_5398_2192.t5 VSS 0.059028f
C1301 a_5398_2192.t0 VSS 0.059028f
C1302 a_5398_2192.n0 VSS 0.139449f
C1303 a_5398_2192.t3 VSS 0.059028f
C1304 a_5398_2192.t1 VSS 0.059028f
C1305 a_5398_2192.n1 VSS 0.258102f
C1306 a_5398_2192.n2 VSS 1.11221f
C1307 a_5398_2192.n3 VSS 0.136068f
C1308 a_5398_2192.t4 VSS 0.059028f
C1309 a_5134_2192.t1 VSS 0.024913f
C1310 a_5134_2192.t5 VSS 0.024913f
C1311 a_5134_2192.t4 VSS 0.024913f
C1312 a_5134_2192.n0 VSS 0.057409f
C1313 a_5134_2192.t6 VSS 0.024913f
C1314 a_5134_2192.t7 VSS 0.024913f
C1315 a_5134_2192.n1 VSS 0.060272f
C1316 a_5134_2192.n2 VSS 0.340434f
C1317 a_5134_2192.t0 VSS 0.024913f
C1318 a_5134_2192.t11 VSS 0.024913f
C1319 a_5134_2192.n3 VSS 0.060114f
C1320 a_5134_2192.t9 VSS 0.024913f
C1321 a_5134_2192.t3 VSS 0.024913f
C1322 a_5134_2192.n4 VSS 0.060114f
C1323 a_5134_2192.t2 VSS 0.024913f
C1324 a_5134_2192.t12 VSS 0.024913f
C1325 a_5134_2192.n5 VSS 0.060114f
C1326 a_5134_2192.t10 VSS 0.097139f
C1327 a_5134_2192.n6 VSS 0.369186f
C1328 a_5134_2192.n7 VSS 0.182473f
C1329 a_5134_2192.n8 VSS 0.22019f
C1330 a_5134_2192.n9 VSS 0.140942f
C1331 a_5134_2192.n10 VSS 0.052659f
C1332 a_5134_2192.t8 VSS 0.024913f
C1333 saff_delay_unit_1/delay_unit_2_0.in_1.t13 VSS 0.060272f
C1334 saff_delay_unit_1/delay_unit_2_0.in_1.t17 VSS 0.018895f
C1335 saff_delay_unit_1/delay_unit_2_0.in_1.n0 VSS 0.044259f
C1336 saff_delay_unit_1/delay_unit_2_0.in_1.t10 VSS 0.060272f
C1337 saff_delay_unit_1/delay_unit_2_0.in_1.t12 VSS 0.018895f
C1338 saff_delay_unit_1/delay_unit_2_0.in_1.n1 VSS 0.044618f
C1339 saff_delay_unit_1/delay_unit_2_0.in_1.n2 VSS 0.017344f
C1340 saff_delay_unit_1/delay_unit_2_0.in_1.t16 VSS 0.060272f
C1341 saff_delay_unit_1/delay_unit_2_0.in_1.t19 VSS 0.018895f
C1342 saff_delay_unit_1/delay_unit_2_0.in_1.n3 VSS 0.044618f
C1343 saff_delay_unit_1/delay_unit_2_0.in_1.t9 VSS 0.060272f
C1344 saff_delay_unit_1/delay_unit_2_0.in_1.t11 VSS 0.018895f
C1345 saff_delay_unit_1/delay_unit_2_0.in_1.n4 VSS 0.044259f
C1346 saff_delay_unit_1/delay_unit_2_0.in_1.n5 VSS 0.017194f
C1347 saff_delay_unit_1/delay_unit_2_0.in_1.n6 VSS 0.355789f
C1348 saff_delay_unit_1/delay_unit_2_0.in_1.t6 VSS 0.048788f
C1349 saff_delay_unit_1/delay_unit_2_0.in_1.t7 VSS 0.147676f
C1350 saff_delay_unit_1/delay_unit_2_0.in_1.n7 VSS 0.374807f
C1351 saff_delay_unit_1/delay_unit_2_0.in_1.n8 VSS 0.193404f
C1352 saff_delay_unit_1/delay_unit_2_0.in_1.t2 VSS 0.013333f
C1353 saff_delay_unit_1/delay_unit_2_0.in_1.t1 VSS 0.013333f
C1354 saff_delay_unit_1/delay_unit_2_0.in_1.n9 VSS 0.031228f
C1355 saff_delay_unit_1/delay_unit_2_0.in_1.t5 VSS 0.039998f
C1356 saff_delay_unit_1/delay_unit_2_0.in_1.t4 VSS 0.039998f
C1357 saff_delay_unit_1/delay_unit_2_0.in_1.n10 VSS 0.081482f
C1358 saff_delay_unit_1/delay_unit_2_0.in_1.n11 VSS 0.339017f
C1359 saff_delay_unit_1/delay_unit_2_0.in_1.t18 VSS 0.062608f
C1360 saff_delay_unit_1/delay_unit_2_0.in_1.t14 VSS 0.062608f
C1361 saff_delay_unit_1/delay_unit_2_0.in_1.n12 VSS 0.070681f
C1362 saff_delay_unit_1/delay_unit_2_0.in_1.t15 VSS 0.062608f
C1363 saff_delay_unit_1/delay_unit_2_0.in_1.t8 VSS 0.062608f
C1364 saff_delay_unit_1/delay_unit_2_0.in_1.n13 VSS 0.070298f
C1365 saff_delay_unit_1/delay_unit_2_0.in_1.n14 VSS 0.641836f
C1366 saff_delay_unit_1/delay_unit_2_0.in_1.t0 VSS 0.046823f
C1367 saff_delay_unit_1/delay_unit_2_0.in_1.n15 VSS 0.161715f
C1368 saff_delay_unit_1/delay_unit_2_0.in_1.t3 VSS 0.147676f
C1369 saff_delay_unit_1/delay_unit_2_0.in_1.n16 VSS 0.245085f
C1370 saff_delay_unit_1/delay_unit_2_0.in_1.n17 VSS 0.184206f
C1371 saff_delay_unit_2/delay_unit_2_0.in_2.t12 VSS 0.039951f
C1372 saff_delay_unit_2/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1373 saff_delay_unit_2/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1374 saff_delay_unit_2/delay_unit_2_0.in_2.t13 VSS 0.039951f
C1375 saff_delay_unit_2/delay_unit_2_0.in_2.t17 VSS 0.012525f
C1376 saff_delay_unit_2/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1377 saff_delay_unit_2/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1378 saff_delay_unit_2/delay_unit_2_0.in_2.t19 VSS 0.039951f
C1379 saff_delay_unit_2/delay_unit_2_0.in_2.t8 VSS 0.012525f
C1380 saff_delay_unit_2/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1381 saff_delay_unit_2/delay_unit_2_0.in_2.t11 VSS 0.039951f
C1382 saff_delay_unit_2/delay_unit_2_0.in_2.t14 VSS 0.012525f
C1383 saff_delay_unit_2/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1384 saff_delay_unit_2/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1385 saff_delay_unit_2/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1386 saff_delay_unit_2/delay_unit_2_0.in_2.t7 VSS 0.100425f
C1387 saff_delay_unit_2/delay_unit_2_0.in_2.t6 VSS 0.031036f
C1388 saff_delay_unit_2/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1389 saff_delay_unit_2/delay_unit_2_0.in_2.t9 VSS 0.047479f
C1390 saff_delay_unit_2/delay_unit_2_0.in_2.t16 VSS 0.047479f
C1391 saff_delay_unit_2/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1392 saff_delay_unit_2/delay_unit_2_0.in_2.t10 VSS 0.047479f
C1393 saff_delay_unit_2/delay_unit_2_0.in_2.t18 VSS 0.047479f
C1394 saff_delay_unit_2/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1395 saff_delay_unit_2/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1396 saff_delay_unit_2/delay_unit_2_0.in_2.t5 VSS 0.026512f
C1397 saff_delay_unit_2/delay_unit_2_0.in_2.t2 VSS 0.026512f
C1398 saff_delay_unit_2/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1399 saff_delay_unit_2/delay_unit_2_0.in_2.t4 VSS 0.008837f
C1400 saff_delay_unit_2/delay_unit_2_0.in_2.t0 VSS 0.008837f
C1401 saff_delay_unit_2/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1402 saff_delay_unit_2/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1403 saff_delay_unit_2/delay_unit_2_0.in_2.t3 VSS 0.100425f
C1404 saff_delay_unit_2/delay_unit_2_0.in_2.t1 VSS 0.031036f
C1405 saff_delay_unit_2/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1406 saff_delay_unit_2/delay_unit_2_0.in_2.n15 VSS 0.126574f
C1407 a_16808_2192.t5 VSS 0.059028f
C1408 a_16808_2192.t2 VSS 0.059028f
C1409 a_16808_2192.t0 VSS 0.059028f
C1410 a_16808_2192.n0 VSS 0.136068f
C1411 a_16808_2192.t3 VSS 0.059028f
C1412 a_16808_2192.t1 VSS 0.059028f
C1413 a_16808_2192.n1 VSS 0.258102f
C1414 a_16808_2192.n2 VSS 1.11221f
C1415 a_16808_2192.n3 VSS 0.139449f
C1416 a_16808_2192.t4 VSS 0.059028f
C1417 saff_delay_unit_3/delay_unit_2_0.in_1.t9 VSS 0.059113f
C1418 saff_delay_unit_3/delay_unit_2_0.in_1.t11 VSS 0.018532f
C1419 saff_delay_unit_3/delay_unit_2_0.in_1.n0 VSS 0.043408f
C1420 saff_delay_unit_3/delay_unit_2_0.in_1.t15 VSS 0.059113f
C1421 saff_delay_unit_3/delay_unit_2_0.in_1.t17 VSS 0.018532f
C1422 saff_delay_unit_3/delay_unit_2_0.in_1.n1 VSS 0.04376f
C1423 saff_delay_unit_3/delay_unit_2_0.in_1.n2 VSS 0.01701f
C1424 saff_delay_unit_3/delay_unit_2_0.in_1.t8 VSS 0.059113f
C1425 saff_delay_unit_3/delay_unit_2_0.in_1.t10 VSS 0.018532f
C1426 saff_delay_unit_3/delay_unit_2_0.in_1.n3 VSS 0.04376f
C1427 saff_delay_unit_3/delay_unit_2_0.in_1.t13 VSS 0.059113f
C1428 saff_delay_unit_3/delay_unit_2_0.in_1.t16 VSS 0.018532f
C1429 saff_delay_unit_3/delay_unit_2_0.in_1.n4 VSS 0.043408f
C1430 saff_delay_unit_3/delay_unit_2_0.in_1.n5 VSS 0.016864f
C1431 saff_delay_unit_3/delay_unit_2_0.in_1.n6 VSS 0.348947f
C1432 saff_delay_unit_3/delay_unit_2_0.in_1.t6 VSS 0.04785f
C1433 saff_delay_unit_3/delay_unit_2_0.in_1.t7 VSS 0.144836f
C1434 saff_delay_unit_3/delay_unit_2_0.in_1.n7 VSS 0.367599f
C1435 saff_delay_unit_3/delay_unit_2_0.in_1.t2 VSS 0.013076f
C1436 saff_delay_unit_3/delay_unit_2_0.in_1.t4 VSS 0.013076f
C1437 saff_delay_unit_3/delay_unit_2_0.in_1.n8 VSS 0.030628f
C1438 saff_delay_unit_3/delay_unit_2_0.in_1.t0 VSS 0.039228f
C1439 saff_delay_unit_3/delay_unit_2_0.in_1.t3 VSS 0.039228f
C1440 saff_delay_unit_3/delay_unit_2_0.in_1.n9 VSS 0.079915f
C1441 saff_delay_unit_3/delay_unit_2_0.in_1.n10 VSS 0.332497f
C1442 saff_delay_unit_3/delay_unit_2_0.in_1.t14 VSS 0.061404f
C1443 saff_delay_unit_3/delay_unit_2_0.in_1.t19 VSS 0.061404f
C1444 saff_delay_unit_3/delay_unit_2_0.in_1.n11 VSS 0.069322f
C1445 saff_delay_unit_3/delay_unit_2_0.in_1.t12 VSS 0.061404f
C1446 saff_delay_unit_3/delay_unit_2_0.in_1.t18 VSS 0.061404f
C1447 saff_delay_unit_3/delay_unit_2_0.in_1.n12 VSS 0.068946f
C1448 saff_delay_unit_3/delay_unit_2_0.in_1.n13 VSS 0.629493f
C1449 saff_delay_unit_3/delay_unit_2_0.in_1.t1 VSS 0.045922f
C1450 saff_delay_unit_3/delay_unit_2_0.in_1.n14 VSS 0.158606f
C1451 saff_delay_unit_3/delay_unit_2_0.in_1.t5 VSS 0.144836f
C1452 saff_delay_unit_3/delay_unit_2_0.in_1.n15 VSS 0.240372f
C1453 saff_delay_unit_3/delay_unit_2_0.in_1.n16 VSS 0.180663f
C1454 saff_delay_unit_5/delay_unit_2_0.in_2.t18 VSS 0.039951f
C1455 saff_delay_unit_5/delay_unit_2_0.in_2.t9 VSS 0.012525f
C1456 saff_delay_unit_5/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1457 saff_delay_unit_5/delay_unit_2_0.in_2.t11 VSS 0.039951f
C1458 saff_delay_unit_5/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1459 saff_delay_unit_5/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1460 saff_delay_unit_5/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1461 saff_delay_unit_5/delay_unit_2_0.in_2.t16 VSS 0.039951f
C1462 saff_delay_unit_5/delay_unit_2_0.in_2.t19 VSS 0.012525f
C1463 saff_delay_unit_5/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1464 saff_delay_unit_5/delay_unit_2_0.in_2.t10 VSS 0.039951f
C1465 saff_delay_unit_5/delay_unit_2_0.in_2.t14 VSS 0.012525f
C1466 saff_delay_unit_5/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1467 saff_delay_unit_5/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1468 saff_delay_unit_5/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1469 saff_delay_unit_5/delay_unit_2_0.in_2.t7 VSS 0.100425f
C1470 saff_delay_unit_5/delay_unit_2_0.in_2.t6 VSS 0.031036f
C1471 saff_delay_unit_5/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1472 saff_delay_unit_5/delay_unit_2_0.in_2.t8 VSS 0.047479f
C1473 saff_delay_unit_5/delay_unit_2_0.in_2.t13 VSS 0.047479f
C1474 saff_delay_unit_5/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1475 saff_delay_unit_5/delay_unit_2_0.in_2.t12 VSS 0.047479f
C1476 saff_delay_unit_5/delay_unit_2_0.in_2.t17 VSS 0.047479f
C1477 saff_delay_unit_5/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1478 saff_delay_unit_5/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1479 saff_delay_unit_5/delay_unit_2_0.in_2.t3 VSS 0.026512f
C1480 saff_delay_unit_5/delay_unit_2_0.in_2.t5 VSS 0.026512f
C1481 saff_delay_unit_5/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1482 saff_delay_unit_5/delay_unit_2_0.in_2.t1 VSS 0.008837f
C1483 saff_delay_unit_5/delay_unit_2_0.in_2.t0 VSS 0.008837f
C1484 saff_delay_unit_5/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1485 saff_delay_unit_5/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1486 saff_delay_unit_5/delay_unit_2_0.in_2.t4 VSS 0.100425f
C1487 saff_delay_unit_5/delay_unit_2_0.in_2.t2 VSS 0.031036f
C1488 saff_delay_unit_5/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1489 saff_delay_unit_5/delay_unit_2_0.in_2.n15 VSS 0.052094f
C1490 saff_delay_unit_5/delay_unit_2_0.in_2.n16 VSS 0.126574f
C1491 saff_delay_unit_4/delay_unit_2_0.in_1.t16 VSS 0.061404f
C1492 saff_delay_unit_4/delay_unit_2_0.in_1.t10 VSS 0.061404f
C1493 saff_delay_unit_4/delay_unit_2_0.in_1.n0 VSS 0.069322f
C1494 saff_delay_unit_4/delay_unit_2_0.in_1.t14 VSS 0.061404f
C1495 saff_delay_unit_4/delay_unit_2_0.in_1.t9 VSS 0.061404f
C1496 saff_delay_unit_4/delay_unit_2_0.in_1.n1 VSS 0.068946f
C1497 saff_delay_unit_4/delay_unit_2_0.in_1.n2 VSS 0.629493f
C1498 saff_delay_unit_4/delay_unit_2_0.in_1.t17 VSS 0.059113f
C1499 saff_delay_unit_4/delay_unit_2_0.in_1.t8 VSS 0.018532f
C1500 saff_delay_unit_4/delay_unit_2_0.in_1.n3 VSS 0.043408f
C1501 saff_delay_unit_4/delay_unit_2_0.in_1.t19 VSS 0.059113f
C1502 saff_delay_unit_4/delay_unit_2_0.in_1.t12 VSS 0.018532f
C1503 saff_delay_unit_4/delay_unit_2_0.in_1.n4 VSS 0.04376f
C1504 saff_delay_unit_4/delay_unit_2_0.in_1.n5 VSS 0.01701f
C1505 saff_delay_unit_4/delay_unit_2_0.in_1.t13 VSS 0.059113f
C1506 saff_delay_unit_4/delay_unit_2_0.in_1.t15 VSS 0.018532f
C1507 saff_delay_unit_4/delay_unit_2_0.in_1.n6 VSS 0.04376f
C1508 saff_delay_unit_4/delay_unit_2_0.in_1.t18 VSS 0.059113f
C1509 saff_delay_unit_4/delay_unit_2_0.in_1.t11 VSS 0.018532f
C1510 saff_delay_unit_4/delay_unit_2_0.in_1.n7 VSS 0.043408f
C1511 saff_delay_unit_4/delay_unit_2_0.in_1.n8 VSS 0.016864f
C1512 saff_delay_unit_4/delay_unit_2_0.in_1.n9 VSS 0.348947f
C1513 saff_delay_unit_4/delay_unit_2_0.in_1.t6 VSS 0.04785f
C1514 saff_delay_unit_4/delay_unit_2_0.in_1.t7 VSS 0.144836f
C1515 saff_delay_unit_4/delay_unit_2_0.in_1.n10 VSS 0.367599f
C1516 saff_delay_unit_4/delay_unit_2_0.in_1.n11 VSS 0.189684f
C1517 saff_delay_unit_4/delay_unit_2_0.in_1.t2 VSS 0.013076f
C1518 saff_delay_unit_4/delay_unit_2_0.in_1.t0 VSS 0.013076f
C1519 saff_delay_unit_4/delay_unit_2_0.in_1.n12 VSS 0.030628f
C1520 saff_delay_unit_4/delay_unit_2_0.in_1.t3 VSS 0.039228f
C1521 saff_delay_unit_4/delay_unit_2_0.in_1.t4 VSS 0.039228f
C1522 saff_delay_unit_4/delay_unit_2_0.in_1.n13 VSS 0.079915f
C1523 saff_delay_unit_4/delay_unit_2_0.in_1.n14 VSS 0.332497f
C1524 saff_delay_unit_4/delay_unit_2_0.in_1.n15 VSS 0.180663f
C1525 saff_delay_unit_4/delay_unit_2_0.in_1.t5 VSS 0.144836f
C1526 saff_delay_unit_4/delay_unit_2_0.in_1.n16 VSS 0.240372f
C1527 saff_delay_unit_4/delay_unit_2_0.in_1.t1 VSS 0.045922f
C1528 saff_delay_unit_4/delay_unit_2_0.in_1.n17 VSS 0.158606f
C1529 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1530 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1531 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.087567f
C1532 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.039891f
C1533 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1534 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1535 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C1536 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C1537 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.115133f
C1538 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.095888f
C1539 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.041221f
C1540 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.116123f
C1541 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.108538f
C1542 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.081767f
C1543 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.090596f
C1544 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.106694f
C1545 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C1546 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1547 a_2852_2192.t5 VSS 0.024913f
C1548 a_2852_2192.t7 VSS 0.024913f
C1549 a_2852_2192.t6 VSS 0.024913f
C1550 a_2852_2192.n0 VSS 0.057409f
C1551 a_2852_2192.t1 VSS 0.024913f
C1552 a_2852_2192.t11 VSS 0.024913f
C1553 a_2852_2192.n1 VSS 0.060114f
C1554 a_2852_2192.t9 VSS 0.024913f
C1555 a_2852_2192.t2 VSS 0.024913f
C1556 a_2852_2192.n2 VSS 0.060114f
C1557 a_2852_2192.t0 VSS 0.024913f
C1558 a_2852_2192.t10 VSS 0.024913f
C1559 a_2852_2192.n3 VSS 0.060114f
C1560 a_2852_2192.t12 VSS 0.097139f
C1561 a_2852_2192.n4 VSS 0.369186f
C1562 a_2852_2192.n5 VSS 0.182473f
C1563 a_2852_2192.n6 VSS 0.22019f
C1564 a_2852_2192.t4 VSS 0.024913f
C1565 a_2852_2192.t3 VSS 0.024913f
C1566 a_2852_2192.n7 VSS 0.052659f
C1567 a_2852_2192.n8 VSS 0.140942f
C1568 a_2852_2192.n9 VSS 0.340434f
C1569 a_2852_2192.n10 VSS 0.060272f
C1570 a_2852_2192.t8 VSS 0.024913f
C1571 a_14262_2192.t8 VSS 0.024913f
C1572 a_14262_2192.t9 VSS 0.024913f
C1573 a_14262_2192.t12 VSS 0.024913f
C1574 a_14262_2192.n0 VSS 0.057409f
C1575 a_14262_2192.t4 VSS 0.024913f
C1576 a_14262_2192.t0 VSS 0.024913f
C1577 a_14262_2192.n1 VSS 0.060114f
C1578 a_14262_2192.t2 VSS 0.024913f
C1579 a_14262_2192.t5 VSS 0.024913f
C1580 a_14262_2192.n2 VSS 0.060114f
C1581 a_14262_2192.t7 VSS 0.024913f
C1582 a_14262_2192.t1 VSS 0.024913f
C1583 a_14262_2192.n3 VSS 0.060114f
C1584 a_14262_2192.t3 VSS 0.097139f
C1585 a_14262_2192.n4 VSS 0.369186f
C1586 a_14262_2192.n5 VSS 0.182473f
C1587 a_14262_2192.n6 VSS 0.22019f
C1588 a_14262_2192.t10 VSS 0.024913f
C1589 a_14262_2192.t6 VSS 0.024913f
C1590 a_14262_2192.n7 VSS 0.052659f
C1591 a_14262_2192.n8 VSS 0.140942f
C1592 a_14262_2192.n9 VSS 0.340434f
C1593 a_14262_2192.n10 VSS 0.060272f
C1594 a_14262_2192.t11 VSS 0.024913f
C1595 saff_delay_unit_7/delay_unit_2_0.in_1.t17 VSS 0.061404f
C1596 saff_delay_unit_7/delay_unit_2_0.in_1.t12 VSS 0.061404f
C1597 saff_delay_unit_7/delay_unit_2_0.in_1.n0 VSS 0.069322f
C1598 saff_delay_unit_7/delay_unit_2_0.in_1.t13 VSS 0.061404f
C1599 saff_delay_unit_7/delay_unit_2_0.in_1.t8 VSS 0.061404f
C1600 saff_delay_unit_7/delay_unit_2_0.in_1.n1 VSS 0.068946f
C1601 saff_delay_unit_7/delay_unit_2_0.in_1.n2 VSS 0.629493f
C1602 saff_delay_unit_7/delay_unit_2_0.in_1.t18 VSS 0.059113f
C1603 saff_delay_unit_7/delay_unit_2_0.in_1.t10 VSS 0.018532f
C1604 saff_delay_unit_7/delay_unit_2_0.in_1.n3 VSS 0.043408f
C1605 saff_delay_unit_7/delay_unit_2_0.in_1.t19 VSS 0.059113f
C1606 saff_delay_unit_7/delay_unit_2_0.in_1.t11 VSS 0.018532f
C1607 saff_delay_unit_7/delay_unit_2_0.in_1.n4 VSS 0.04376f
C1608 saff_delay_unit_7/delay_unit_2_0.in_1.n5 VSS 0.01701f
C1609 saff_delay_unit_7/delay_unit_2_0.in_1.t14 VSS 0.059113f
C1610 saff_delay_unit_7/delay_unit_2_0.in_1.t15 VSS 0.018532f
C1611 saff_delay_unit_7/delay_unit_2_0.in_1.n6 VSS 0.04376f
C1612 saff_delay_unit_7/delay_unit_2_0.in_1.t16 VSS 0.059113f
C1613 saff_delay_unit_7/delay_unit_2_0.in_1.t9 VSS 0.018532f
C1614 saff_delay_unit_7/delay_unit_2_0.in_1.n7 VSS 0.043408f
C1615 saff_delay_unit_7/delay_unit_2_0.in_1.n8 VSS 0.016864f
C1616 saff_delay_unit_7/delay_unit_2_0.in_1.n9 VSS 0.348947f
C1617 saff_delay_unit_7/delay_unit_2_0.in_1.t1 VSS 0.04785f
C1618 saff_delay_unit_7/delay_unit_2_0.in_1.t4 VSS 0.144836f
C1619 saff_delay_unit_7/delay_unit_2_0.in_1.n10 VSS 0.367599f
C1620 saff_delay_unit_7/delay_unit_2_0.in_1.t0 VSS 0.013076f
C1621 saff_delay_unit_7/delay_unit_2_0.in_1.t7 VSS 0.013076f
C1622 saff_delay_unit_7/delay_unit_2_0.in_1.n11 VSS 0.030628f
C1623 saff_delay_unit_7/delay_unit_2_0.in_1.t3 VSS 0.039228f
C1624 saff_delay_unit_7/delay_unit_2_0.in_1.t6 VSS 0.039228f
C1625 saff_delay_unit_7/delay_unit_2_0.in_1.n12 VSS 0.079915f
C1626 saff_delay_unit_7/delay_unit_2_0.in_1.n13 VSS 0.332497f
C1627 saff_delay_unit_7/delay_unit_2_0.in_1.n14 VSS 0.180663f
C1628 saff_delay_unit_7/delay_unit_2_0.in_1.t2 VSS 0.144836f
C1629 saff_delay_unit_7/delay_unit_2_0.in_1.n15 VSS 0.240372f
C1630 saff_delay_unit_7/delay_unit_2_0.in_1.t5 VSS 0.045922f
C1631 saff_delay_unit_7/delay_unit_2_0.in_1.n16 VSS 0.158606f
C1632 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1633 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1634 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.087567f
C1635 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.039891f
C1636 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1637 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C1638 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.054262f
C1639 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.115133f
C1640 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.201734f
C1641 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.095888f
C1642 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.041221f
C1643 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.116123f
C1644 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.108538f
C1645 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.081767f
C1646 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.090596f
C1647 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.106694f
C1648 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C1649 saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1650 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C1651 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.087824f
C1652 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.040008f
C1653 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C1654 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.200111f
C1655 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.202807f
C1656 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.096169f
C1657 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.041341f
C1658 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C1659 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.082007f
C1660 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.090862f
C1661 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C1662 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C1663 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.107599f
C1664 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C1665 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C1666 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.054421f
C1667 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C1668 saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
C1669 a_16544_2192.t5 VSS 0.024913f
C1670 a_16544_2192.t7 VSS 0.024913f
C1671 a_16544_2192.t6 VSS 0.024913f
C1672 a_16544_2192.n0 VSS 0.057409f
C1673 a_16544_2192.t0 VSS 0.024913f
C1674 a_16544_2192.t10 VSS 0.024913f
C1675 a_16544_2192.n1 VSS 0.060114f
C1676 a_16544_2192.t9 VSS 0.024913f
C1677 a_16544_2192.t3 VSS 0.024913f
C1678 a_16544_2192.n2 VSS 0.060114f
C1679 a_16544_2192.t1 VSS 0.024913f
C1680 a_16544_2192.t12 VSS 0.024913f
C1681 a_16544_2192.n3 VSS 0.060114f
C1682 a_16544_2192.t11 VSS 0.097139f
C1683 a_16544_2192.n4 VSS 0.369186f
C1684 a_16544_2192.n5 VSS 0.182473f
C1685 a_16544_2192.n6 VSS 0.22019f
C1686 a_16544_2192.t4 VSS 0.024913f
C1687 a_16544_2192.t2 VSS 0.024913f
C1688 a_16544_2192.n7 VSS 0.052659f
C1689 a_16544_2192.n8 VSS 0.140942f
C1690 a_16544_2192.n9 VSS 0.340434f
C1691 a_16544_2192.n10 VSS 0.060272f
C1692 a_16544_2192.t8 VSS 0.024913f
C1693 delay_unit_2_0.in_1 VSS 0.373508f
C1694 saff_delay_unit_7/saff_2_0.sense_amplifier_0.d VSS 0.695927f
C1695 saff_delay_unit_7/saff_2_0.d.t9 VSS 0.059113f
C1696 saff_delay_unit_7/saff_2_0.d.t12 VSS 0.018532f
C1697 saff_delay_unit_7/saff_2_0.d.n0 VSS 0.043408f
C1698 saff_delay_unit_7/saff_2_0.d.t16 VSS 0.059113f
C1699 saff_delay_unit_7/saff_2_0.d.t18 VSS 0.018532f
C1700 saff_delay_unit_7/saff_2_0.d.n1 VSS 0.04376f
C1701 saff_delay_unit_7/saff_2_0.d.n2 VSS 0.01701f
C1702 saff_delay_unit_7/saff_2_0.d.t19 VSS 0.059113f
C1703 saff_delay_unit_7/saff_2_0.d.t11 VSS 0.018532f
C1704 saff_delay_unit_7/saff_2_0.d.n3 VSS 0.04376f
C1705 saff_delay_unit_7/saff_2_0.d.t13 VSS 0.059113f
C1706 saff_delay_unit_7/saff_2_0.d.t17 VSS 0.018532f
C1707 saff_delay_unit_7/saff_2_0.d.n4 VSS 0.043408f
C1708 saff_delay_unit_7/saff_2_0.d.n5 VSS 0.016864f
C1709 saff_delay_unit_7/saff_2_0.d.n6 VSS 0.348947f
C1710 saff_delay_unit_7/saff_2_0.d.t0 VSS 0.04785f
C1711 saff_delay_unit_7/saff_2_0.d.t2 VSS 0.144836f
C1712 saff_delay_unit_7/saff_2_0.d.n7 VSS 0.367599f
C1713 saff_delay_unit_7/saff_2_0.d.t7 VSS 0.013076f
C1714 saff_delay_unit_7/saff_2_0.d.t4 VSS 0.013076f
C1715 saff_delay_unit_7/saff_2_0.d.n8 VSS 0.030628f
C1716 saff_delay_unit_7/saff_2_0.d.t5 VSS 0.039228f
C1717 saff_delay_unit_7/saff_2_0.d.t1 VSS 0.039228f
C1718 saff_delay_unit_7/saff_2_0.d.n9 VSS 0.079915f
C1719 saff_delay_unit_7/saff_2_0.d.n10 VSS 0.332497f
C1720 saff_delay_unit_7/saff_2_0.d.t14 VSS 0.061404f
C1721 saff_delay_unit_7/saff_2_0.d.t15 VSS 0.061404f
C1722 saff_delay_unit_7/saff_2_0.d.n11 VSS 0.069322f
C1723 saff_delay_unit_7/saff_2_0.d.t8 VSS 0.061404f
C1724 saff_delay_unit_7/saff_2_0.d.t10 VSS 0.061404f
C1725 saff_delay_unit_7/saff_2_0.d.n12 VSS 0.068946f
C1726 saff_delay_unit_7/saff_2_0.d.n13 VSS 0.629493f
C1727 saff_delay_unit_7/saff_2_0.d.t3 VSS 0.045922f
C1728 saff_delay_unit_7/saff_2_0.d.n14 VSS 0.158606f
C1729 saff_delay_unit_7/saff_2_0.d.t6 VSS 0.144836f
C1730 saff_delay_unit_7/saff_2_0.d.n15 VSS 0.240372f
C1731 saff_delay_unit_7/saff_2_0.d.n16 VSS 0.180663f
C1732 saff_delay_unit_7/delay_unit_2_0.out_1 VSS 0.271115f
C1733 a_570_2192.t6 VSS 0.024913f
C1734 a_570_2192.t4 VSS 0.024913f
C1735 a_570_2192.t7 VSS 0.024913f
C1736 a_570_2192.n0 VSS 0.060272f
C1737 a_570_2192.t9 VSS 0.024913f
C1738 a_570_2192.t0 VSS 0.024913f
C1739 a_570_2192.n1 VSS 0.060114f
C1740 a_570_2192.t3 VSS 0.024913f
C1741 a_570_2192.t11 VSS 0.024913f
C1742 a_570_2192.n2 VSS 0.060114f
C1743 a_570_2192.t10 VSS 0.024913f
C1744 a_570_2192.t1 VSS 0.024913f
C1745 a_570_2192.n3 VSS 0.060114f
C1746 a_570_2192.t2 VSS 0.097139f
C1747 a_570_2192.n4 VSS 0.369186f
C1748 a_570_2192.n5 VSS 0.182473f
C1749 a_570_2192.n6 VSS 0.22019f
C1750 a_570_2192.t5 VSS 0.024913f
C1751 a_570_2192.t12 VSS 0.024913f
C1752 a_570_2192.n7 VSS 0.052659f
C1753 a_570_2192.n8 VSS 0.140942f
C1754 a_570_2192.n9 VSS 0.340434f
C1755 a_570_2192.n10 VSS 0.057409f
C1756 a_570_2192.t8 VSS 0.024913f
C1757 a_834_2192.t1 VSS 0.059028f
C1758 a_834_2192.t5 VSS 0.059028f
C1759 a_834_2192.t2 VSS 0.059028f
C1760 a_834_2192.n0 VSS 0.136068f
C1761 a_834_2192.t4 VSS 0.059028f
C1762 a_834_2192.t3 VSS 0.059028f
C1763 a_834_2192.n1 VSS 0.258102f
C1764 a_834_2192.n2 VSS 1.11221f
C1765 a_834_2192.n3 VSS 0.139449f
C1766 a_834_2192.t0 VSS 0.059028f
C1767 saff_delay_unit_1/delay_unit_2_0.in_2.t17 VSS 0.039951f
C1768 saff_delay_unit_1/delay_unit_2_0.in_2.t8 VSS 0.012525f
C1769 saff_delay_unit_1/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1770 saff_delay_unit_1/delay_unit_2_0.in_2.t19 VSS 0.039951f
C1771 saff_delay_unit_1/delay_unit_2_0.in_2.t12 VSS 0.012525f
C1772 saff_delay_unit_1/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1773 saff_delay_unit_1/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1774 saff_delay_unit_1/delay_unit_2_0.in_2.t14 VSS 0.039951f
C1775 saff_delay_unit_1/delay_unit_2_0.in_2.t16 VSS 0.012525f
C1776 saff_delay_unit_1/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1777 saff_delay_unit_1/delay_unit_2_0.in_2.t18 VSS 0.039951f
C1778 saff_delay_unit_1/delay_unit_2_0.in_2.t11 VSS 0.012525f
C1779 saff_delay_unit_1/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1780 saff_delay_unit_1/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1781 saff_delay_unit_1/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1782 saff_delay_unit_1/delay_unit_2_0.in_2.t1 VSS 0.100425f
C1783 saff_delay_unit_1/delay_unit_2_0.in_2.t0 VSS 0.031036f
C1784 saff_delay_unit_1/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1785 saff_delay_unit_1/delay_unit_2_0.in_2.t10 VSS 0.047479f
C1786 saff_delay_unit_1/delay_unit_2_0.in_2.t13 VSS 0.047479f
C1787 saff_delay_unit_1/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1788 saff_delay_unit_1/delay_unit_2_0.in_2.t9 VSS 0.047479f
C1789 saff_delay_unit_1/delay_unit_2_0.in_2.t15 VSS 0.047479f
C1790 saff_delay_unit_1/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1791 saff_delay_unit_1/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1792 saff_delay_unit_1/delay_unit_2_0.in_2.t5 VSS 0.026512f
C1793 saff_delay_unit_1/delay_unit_2_0.in_2.t6 VSS 0.026512f
C1794 saff_delay_unit_1/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1795 saff_delay_unit_1/delay_unit_2_0.in_2.t4 VSS 0.008837f
C1796 saff_delay_unit_1/delay_unit_2_0.in_2.t2 VSS 0.008837f
C1797 saff_delay_unit_1/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1798 saff_delay_unit_1/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1799 saff_delay_unit_1/delay_unit_2_0.in_2.t7 VSS 0.100425f
C1800 saff_delay_unit_1/delay_unit_2_0.in_2.t3 VSS 0.031036f
C1801 saff_delay_unit_1/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1802 saff_delay_unit_1/delay_unit_2_0.in_2.n15 VSS 0.052094f
C1803 saff_delay_unit_1/delay_unit_2_0.in_2.n16 VSS 0.126574f
C1804 start_pos.t4 VSS 0.0785f
C1805 start_pos.t6 VSS 0.02461f
C1806 start_pos.n0 VSS 0.057645f
C1807 start_pos.t9 VSS 0.0785f
C1808 start_pos.t3 VSS 0.02461f
C1809 start_pos.n1 VSS 0.058112f
C1810 start_pos.n2 VSS 0.022589f
C1811 start_pos.t5 VSS 0.0785f
C1812 start_pos.t8 VSS 0.02461f
C1813 start_pos.n3 VSS 0.058112f
C1814 start_pos.t7 VSS 0.0785f
C1815 start_pos.t2 VSS 0.02461f
C1816 start_pos.n4 VSS 0.057645f
C1817 start_pos.n5 VSS 0.022394f
C1818 start_pos.n6 VSS 0.463391f
C1819 start_pos.t1 VSS 0.063543f
C1820 start_pos.t0 VSS 0.192338f
C1821 start_pos.n7 VSS 0.48816f
C1822 start_pos.n8 VSS 0.251895f
C1823 saff_delay_unit_3/delay_unit_2_0.in_2.t13 VSS 0.039951f
C1824 saff_delay_unit_3/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1825 saff_delay_unit_3/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1826 saff_delay_unit_3/delay_unit_2_0.in_2.t18 VSS 0.039951f
C1827 saff_delay_unit_3/delay_unit_2_0.in_2.t9 VSS 0.012525f
C1828 saff_delay_unit_3/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1829 saff_delay_unit_3/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1830 saff_delay_unit_3/delay_unit_2_0.in_2.t14 VSS 0.039951f
C1831 saff_delay_unit_3/delay_unit_2_0.in_2.t17 VSS 0.012525f
C1832 saff_delay_unit_3/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1833 saff_delay_unit_3/delay_unit_2_0.in_2.t19 VSS 0.039951f
C1834 saff_delay_unit_3/delay_unit_2_0.in_2.t10 VSS 0.012525f
C1835 saff_delay_unit_3/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1836 saff_delay_unit_3/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1837 saff_delay_unit_3/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1838 saff_delay_unit_3/delay_unit_2_0.in_2.t6 VSS 0.100425f
C1839 saff_delay_unit_3/delay_unit_2_0.in_2.t7 VSS 0.031036f
C1840 saff_delay_unit_3/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1841 saff_delay_unit_3/delay_unit_2_0.in_2.t11 VSS 0.047479f
C1842 saff_delay_unit_3/delay_unit_2_0.in_2.t16 VSS 0.047479f
C1843 saff_delay_unit_3/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1844 saff_delay_unit_3/delay_unit_2_0.in_2.t12 VSS 0.047479f
C1845 saff_delay_unit_3/delay_unit_2_0.in_2.t8 VSS 0.047479f
C1846 saff_delay_unit_3/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1847 saff_delay_unit_3/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1848 saff_delay_unit_3/delay_unit_2_0.in_2.t4 VSS 0.026512f
C1849 saff_delay_unit_3/delay_unit_2_0.in_2.t3 VSS 0.026512f
C1850 saff_delay_unit_3/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1851 saff_delay_unit_3/delay_unit_2_0.in_2.t0 VSS 0.008837f
C1852 saff_delay_unit_3/delay_unit_2_0.in_2.t2 VSS 0.008837f
C1853 saff_delay_unit_3/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1854 saff_delay_unit_3/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1855 saff_delay_unit_3/delay_unit_2_0.in_2.t5 VSS 0.100425f
C1856 saff_delay_unit_3/delay_unit_2_0.in_2.t1 VSS 0.031036f
C1857 saff_delay_unit_3/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1858 saff_delay_unit_3/delay_unit_2_0.in_2.n15 VSS 0.052094f
C1859 saff_delay_unit_3/delay_unit_2_0.in_2.n16 VSS 0.126574f
C1860 saff_delay_unit_2/delay_unit_2_0.in_1.t8 VSS 0.059113f
C1861 saff_delay_unit_2/delay_unit_2_0.in_1.t11 VSS 0.018532f
C1862 saff_delay_unit_2/delay_unit_2_0.in_1.n0 VSS 0.043408f
C1863 saff_delay_unit_2/delay_unit_2_0.in_1.t14 VSS 0.059113f
C1864 saff_delay_unit_2/delay_unit_2_0.in_1.t17 VSS 0.018532f
C1865 saff_delay_unit_2/delay_unit_2_0.in_1.n1 VSS 0.04376f
C1866 saff_delay_unit_2/delay_unit_2_0.in_1.n2 VSS 0.01701f
C1867 saff_delay_unit_2/delay_unit_2_0.in_1.t19 VSS 0.059113f
C1868 saff_delay_unit_2/delay_unit_2_0.in_1.t10 VSS 0.018532f
C1869 saff_delay_unit_2/delay_unit_2_0.in_1.n3 VSS 0.04376f
C1870 saff_delay_unit_2/delay_unit_2_0.in_1.t12 VSS 0.059113f
C1871 saff_delay_unit_2/delay_unit_2_0.in_1.t15 VSS 0.018532f
C1872 saff_delay_unit_2/delay_unit_2_0.in_1.n4 VSS 0.043408f
C1873 saff_delay_unit_2/delay_unit_2_0.in_1.n5 VSS 0.016864f
C1874 saff_delay_unit_2/delay_unit_2_0.in_1.n6 VSS 0.348947f
C1875 saff_delay_unit_2/delay_unit_2_0.in_1.t0 VSS 0.04785f
C1876 saff_delay_unit_2/delay_unit_2_0.in_1.t1 VSS 0.144836f
C1877 saff_delay_unit_2/delay_unit_2_0.in_1.n7 VSS 0.367599f
C1878 saff_delay_unit_2/delay_unit_2_0.in_1.t6 VSS 0.013076f
C1879 saff_delay_unit_2/delay_unit_2_0.in_1.t2 VSS 0.013076f
C1880 saff_delay_unit_2/delay_unit_2_0.in_1.n8 VSS 0.030628f
C1881 saff_delay_unit_2/delay_unit_2_0.in_1.t3 VSS 0.039228f
C1882 saff_delay_unit_2/delay_unit_2_0.in_1.t7 VSS 0.039228f
C1883 saff_delay_unit_2/delay_unit_2_0.in_1.n9 VSS 0.079915f
C1884 saff_delay_unit_2/delay_unit_2_0.in_1.n10 VSS 0.332497f
C1885 saff_delay_unit_2/delay_unit_2_0.in_1.t13 VSS 0.061404f
C1886 saff_delay_unit_2/delay_unit_2_0.in_1.t18 VSS 0.061404f
C1887 saff_delay_unit_2/delay_unit_2_0.in_1.n11 VSS 0.069322f
C1888 saff_delay_unit_2/delay_unit_2_0.in_1.t16 VSS 0.061404f
C1889 saff_delay_unit_2/delay_unit_2_0.in_1.t9 VSS 0.061404f
C1890 saff_delay_unit_2/delay_unit_2_0.in_1.n12 VSS 0.068946f
C1891 saff_delay_unit_2/delay_unit_2_0.in_1.n13 VSS 0.629493f
C1892 saff_delay_unit_2/delay_unit_2_0.in_1.t5 VSS 0.045922f
C1893 saff_delay_unit_2/delay_unit_2_0.in_1.n14 VSS 0.158606f
C1894 saff_delay_unit_2/delay_unit_2_0.in_1.t4 VSS 0.144836f
C1895 saff_delay_unit_2/delay_unit_2_0.in_1.n15 VSS 0.240372f
C1896 saff_delay_unit_2/delay_unit_2_0.in_1.n16 VSS 0.180663f
C1897 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1898 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1899 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.087567f
C1900 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.039891f
C1901 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1902 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1903 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C1904 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.095888f
C1905 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.041221f
C1906 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C1907 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.108538f
C1908 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.081767f
C1909 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.090596f
C1910 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C1911 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C1912 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C1913 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C1914 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1915 saff_delay_unit_5/delay_unit_2_0.in_1.t19 VSS 0.059113f
C1916 saff_delay_unit_5/delay_unit_2_0.in_1.t9 VSS 0.018532f
C1917 saff_delay_unit_5/delay_unit_2_0.in_1.n0 VSS 0.043408f
C1918 saff_delay_unit_5/delay_unit_2_0.in_1.t13 VSS 0.059113f
C1919 saff_delay_unit_5/delay_unit_2_0.in_1.t16 VSS 0.018532f
C1920 saff_delay_unit_5/delay_unit_2_0.in_1.n1 VSS 0.04376f
C1921 saff_delay_unit_5/delay_unit_2_0.in_1.n2 VSS 0.01701f
C1922 saff_delay_unit_5/delay_unit_2_0.in_1.t17 VSS 0.059113f
C1923 saff_delay_unit_5/delay_unit_2_0.in_1.t8 VSS 0.018532f
C1924 saff_delay_unit_5/delay_unit_2_0.in_1.n3 VSS 0.04376f
C1925 saff_delay_unit_5/delay_unit_2_0.in_1.t11 VSS 0.059113f
C1926 saff_delay_unit_5/delay_unit_2_0.in_1.t15 VSS 0.018532f
C1927 saff_delay_unit_5/delay_unit_2_0.in_1.n4 VSS 0.043408f
C1928 saff_delay_unit_5/delay_unit_2_0.in_1.n5 VSS 0.016864f
C1929 saff_delay_unit_5/delay_unit_2_0.in_1.n6 VSS 0.348947f
C1930 saff_delay_unit_5/delay_unit_2_0.in_1.t0 VSS 0.04785f
C1931 saff_delay_unit_5/delay_unit_2_0.in_1.t7 VSS 0.144836f
C1932 saff_delay_unit_5/delay_unit_2_0.in_1.n7 VSS 0.367599f
C1933 saff_delay_unit_5/delay_unit_2_0.in_1.n8 VSS 0.189684f
C1934 saff_delay_unit_5/delay_unit_2_0.in_1.t2 VSS 0.013076f
C1935 saff_delay_unit_5/delay_unit_2_0.in_1.t3 VSS 0.013076f
C1936 saff_delay_unit_5/delay_unit_2_0.in_1.n9 VSS 0.030628f
C1937 saff_delay_unit_5/delay_unit_2_0.in_1.t6 VSS 0.039228f
C1938 saff_delay_unit_5/delay_unit_2_0.in_1.t4 VSS 0.039228f
C1939 saff_delay_unit_5/delay_unit_2_0.in_1.n10 VSS 0.079915f
C1940 saff_delay_unit_5/delay_unit_2_0.in_1.n11 VSS 0.332497f
C1941 saff_delay_unit_5/delay_unit_2_0.in_1.t10 VSS 0.061404f
C1942 saff_delay_unit_5/delay_unit_2_0.in_1.t14 VSS 0.061404f
C1943 saff_delay_unit_5/delay_unit_2_0.in_1.n12 VSS 0.069322f
C1944 saff_delay_unit_5/delay_unit_2_0.in_1.t18 VSS 0.061404f
C1945 saff_delay_unit_5/delay_unit_2_0.in_1.t12 VSS 0.061404f
C1946 saff_delay_unit_5/delay_unit_2_0.in_1.n13 VSS 0.068946f
C1947 saff_delay_unit_5/delay_unit_2_0.in_1.n14 VSS 0.629493f
C1948 saff_delay_unit_5/delay_unit_2_0.in_1.t1 VSS 0.045922f
C1949 saff_delay_unit_5/delay_unit_2_0.in_1.n15 VSS 0.158606f
C1950 saff_delay_unit_5/delay_unit_2_0.in_1.t5 VSS 0.144836f
C1951 saff_delay_unit_5/delay_unit_2_0.in_1.n16 VSS 0.240372f
C1952 saff_delay_unit_5/delay_unit_2_0.in_1.n17 VSS 0.180663f
C1953 saff_delay_unit_4/delay_unit_2_0.in_2.t17 VSS 0.039951f
C1954 saff_delay_unit_4/delay_unit_2_0.in_2.t19 VSS 0.012525f
C1955 saff_delay_unit_4/delay_unit_2_0.in_2.n0 VSS 0.029574f
C1956 saff_delay_unit_4/delay_unit_2_0.in_2.t11 VSS 0.039951f
C1957 saff_delay_unit_4/delay_unit_2_0.in_2.t15 VSS 0.012525f
C1958 saff_delay_unit_4/delay_unit_2_0.in_2.n1 VSS 0.029337f
C1959 saff_delay_unit_4/delay_unit_2_0.in_2.n2 VSS 0.011494f
C1960 saff_delay_unit_4/delay_unit_2_0.in_2.t18 VSS 0.039951f
C1961 saff_delay_unit_4/delay_unit_2_0.in_2.t8 VSS 0.012525f
C1962 saff_delay_unit_4/delay_unit_2_0.in_2.n3 VSS 0.029574f
C1963 saff_delay_unit_4/delay_unit_2_0.in_2.t9 VSS 0.039951f
C1964 saff_delay_unit_4/delay_unit_2_0.in_2.t13 VSS 0.012525f
C1965 saff_delay_unit_4/delay_unit_2_0.in_2.n4 VSS 0.029337f
C1966 saff_delay_unit_4/delay_unit_2_0.in_2.n5 VSS 0.011397f
C1967 saff_delay_unit_4/delay_unit_2_0.in_2.n6 VSS 0.138751f
C1968 saff_delay_unit_4/delay_unit_2_0.in_2.t7 VSS 0.100425f
C1969 saff_delay_unit_4/delay_unit_2_0.in_2.t6 VSS 0.031036f
C1970 saff_delay_unit_4/delay_unit_2_0.in_2.n7 VSS 0.274483f
C1971 saff_delay_unit_4/delay_unit_2_0.in_2.t14 VSS 0.047479f
C1972 saff_delay_unit_4/delay_unit_2_0.in_2.t10 VSS 0.047479f
C1973 saff_delay_unit_4/delay_unit_2_0.in_2.n8 VSS 0.055625f
C1974 saff_delay_unit_4/delay_unit_2_0.in_2.t12 VSS 0.047479f
C1975 saff_delay_unit_4/delay_unit_2_0.in_2.t16 VSS 0.047479f
C1976 saff_delay_unit_4/delay_unit_2_0.in_2.n9 VSS 0.055374f
C1977 saff_delay_unit_4/delay_unit_2_0.in_2.n10 VSS 0.507513f
C1978 saff_delay_unit_4/delay_unit_2_0.in_2.t3 VSS 0.026512f
C1979 saff_delay_unit_4/delay_unit_2_0.in_2.t5 VSS 0.026512f
C1980 saff_delay_unit_4/delay_unit_2_0.in_2.n11 VSS 0.056695f
C1981 saff_delay_unit_4/delay_unit_2_0.in_2.t1 VSS 0.008837f
C1982 saff_delay_unit_4/delay_unit_2_0.in_2.t2 VSS 0.008837f
C1983 saff_delay_unit_4/delay_unit_2_0.in_2.n12 VSS 0.019186f
C1984 saff_delay_unit_4/delay_unit_2_0.in_2.n13 VSS 0.227994f
C1985 saff_delay_unit_4/delay_unit_2_0.in_2.t0 VSS 0.100425f
C1986 saff_delay_unit_4/delay_unit_2_0.in_2.t4 VSS 0.031036f
C1987 saff_delay_unit_4/delay_unit_2_0.in_2.n14 VSS 0.241348f
C1988 saff_delay_unit_4/delay_unit_2_0.in_2.n15 VSS 0.126574f
C1989 a_11980_2192.t8 VSS 0.024913f
C1990 a_11980_2192.t7 VSS 0.024913f
C1991 a_11980_2192.t6 VSS 0.024913f
C1992 a_11980_2192.n0 VSS 0.060272f
C1993 a_11980_2192.t12 VSS 0.024913f
C1994 a_11980_2192.t5 VSS 0.024913f
C1995 a_11980_2192.n1 VSS 0.060114f
C1996 a_11980_2192.t4 VSS 0.024913f
C1997 a_11980_2192.t1 VSS 0.024913f
C1998 a_11980_2192.n2 VSS 0.060114f
C1999 a_11980_2192.t3 VSS 0.024913f
C2000 a_11980_2192.t2 VSS 0.024913f
C2001 a_11980_2192.n3 VSS 0.060114f
C2002 a_11980_2192.t0 VSS 0.097139f
C2003 a_11980_2192.n4 VSS 0.369186f
C2004 a_11980_2192.n5 VSS 0.182473f
C2005 a_11980_2192.n6 VSS 0.22019f
C2006 a_11980_2192.t9 VSS 0.024913f
C2007 a_11980_2192.t11 VSS 0.024913f
C2008 a_11980_2192.n7 VSS 0.052659f
C2009 a_11980_2192.n8 VSS 0.140942f
C2010 a_11980_2192.n9 VSS 0.340434f
C2011 a_11980_2192.n10 VSS 0.057409f
C2012 a_11980_2192.t10 VSS 0.024913f
C2013 stop_strong.t25 VSS 0.075034f
C2014 stop_strong.t27 VSS 0.074865f
C2015 stop_strong.n0 VSS 0.322903f
C2016 stop_strong.t2 VSS 0.057644f
C2017 stop_strong.t42 VSS 0.057644f
C2018 stop_strong.t8 VSS 0.057644f
C2019 stop_strong.t32 VSS 0.057644f
C2020 stop_strong.t44 VSS 0.063869f
C2021 stop_strong.n1 VSS 0.056168f
C2022 stop_strong.n2 VSS 0.033109f
C2023 stop_strong.n3 VSS 0.033109f
C2024 stop_strong.n4 VSS 0.049874f
C2025 stop_strong.n5 VSS 0.749968f
C2026 stop_strong.t15 VSS 0.075034f
C2027 stop_strong.t55 VSS 0.074865f
C2028 stop_strong.n6 VSS 0.322903f
C2029 stop_strong.t50 VSS 0.057644f
C2030 stop_strong.t17 VSS 0.057644f
C2031 stop_strong.t43 VSS 0.057644f
C2032 stop_strong.t9 VSS 0.057644f
C2033 stop_strong.t33 VSS 0.063869f
C2034 stop_strong.n7 VSS 0.056168f
C2035 stop_strong.n8 VSS 0.033109f
C2036 stop_strong.n9 VSS 0.033109f
C2037 stop_strong.n10 VSS 0.049874f
C2038 stop_strong.n11 VSS 0.625244f
C2039 stop_strong.n12 VSS 0.558556f
C2040 stop_strong.t49 VSS 0.075034f
C2041 stop_strong.t45 VSS 0.074865f
C2042 stop_strong.n13 VSS 0.322903f
C2043 stop_strong.t39 VSS 0.057644f
C2044 stop_strong.t51 VSS 0.057644f
C2045 stop_strong.t0 VSS 0.057644f
C2046 stop_strong.t37 VSS 0.057644f
C2047 stop_strong.t3 VSS 0.063869f
C2048 stop_strong.n14 VSS 0.056168f
C2049 stop_strong.n15 VSS 0.033109f
C2050 stop_strong.n16 VSS 0.033109f
C2051 stop_strong.n17 VSS 0.049874f
C2052 stop_strong.n18 VSS 0.625244f
C2053 stop_strong.n19 VSS 0.558556f
C2054 stop_strong.t28 VSS 0.075034f
C2055 stop_strong.t34 VSS 0.074865f
C2056 stop_strong.n20 VSS 0.322903f
C2057 stop_strong.t53 VSS 0.057644f
C2058 stop_strong.t20 VSS 0.057644f
C2059 stop_strong.t46 VSS 0.057644f
C2060 stop_strong.t11 VSS 0.057644f
C2061 stop_strong.t52 VSS 0.063869f
C2062 stop_strong.n21 VSS 0.056168f
C2063 stop_strong.n22 VSS 0.033109f
C2064 stop_strong.n23 VSS 0.033109f
C2065 stop_strong.n24 VSS 0.049874f
C2066 stop_strong.n25 VSS 0.625244f
C2067 stop_strong.n26 VSS 0.558556f
C2068 stop_strong.t19 VSS 0.075034f
C2069 stop_strong.t35 VSS 0.074865f
C2070 stop_strong.n27 VSS 0.322903f
C2071 stop_strong.t54 VSS 0.057644f
C2072 stop_strong.t21 VSS 0.057644f
C2073 stop_strong.t47 VSS 0.057644f
C2074 stop_strong.t12 VSS 0.057644f
C2075 stop_strong.t38 VSS 0.063869f
C2076 stop_strong.n28 VSS 0.056168f
C2077 stop_strong.n29 VSS 0.033109f
C2078 stop_strong.n30 VSS 0.033109f
C2079 stop_strong.n31 VSS 0.049874f
C2080 stop_strong.n32 VSS 0.625244f
C2081 stop_strong.n33 VSS 0.558556f
C2082 stop_strong.t6 VSS 0.075034f
C2083 stop_strong.t31 VSS 0.074865f
C2084 stop_strong.n34 VSS 0.322903f
C2085 stop_strong.t29 VSS 0.057644f
C2086 stop_strong.t10 VSS 0.057644f
C2087 stop_strong.t36 VSS 0.057644f
C2088 stop_strong.t40 VSS 0.057644f
C2089 stop_strong.t7 VSS 0.063869f
C2090 stop_strong.n35 VSS 0.056168f
C2091 stop_strong.n36 VSS 0.033109f
C2092 stop_strong.n37 VSS 0.033109f
C2093 stop_strong.n38 VSS 0.049874f
C2094 stop_strong.n39 VSS 0.625244f
C2095 stop_strong.n40 VSS 0.558556f
C2096 stop_strong.t22 VSS 0.075034f
C2097 stop_strong.t23 VSS 0.074865f
C2098 stop_strong.n41 VSS 0.322903f
C2099 stop_strong.t1 VSS 0.057644f
C2100 stop_strong.t24 VSS 0.057644f
C2101 stop_strong.t4 VSS 0.057644f
C2102 stop_strong.t16 VSS 0.057644f
C2103 stop_strong.t41 VSS 0.063869f
C2104 stop_strong.n42 VSS 0.056168f
C2105 stop_strong.n43 VSS 0.033109f
C2106 stop_strong.n44 VSS 0.033109f
C2107 stop_strong.n45 VSS 0.049874f
C2108 stop_strong.n46 VSS 0.625244f
C2109 stop_strong.n47 VSS 0.558556f
C2110 stop_strong.t18 VSS 0.075034f
C2111 stop_strong.t13 VSS 0.074865f
C2112 stop_strong.n48 VSS 0.322903f
C2113 stop_strong.t48 VSS 0.057644f
C2114 stop_strong.t14 VSS 0.057644f
C2115 stop_strong.t26 VSS 0.057644f
C2116 stop_strong.t5 VSS 0.057644f
C2117 stop_strong.t30 VSS 0.063869f
C2118 stop_strong.n49 VSS 0.056168f
C2119 stop_strong.n50 VSS 0.033109f
C2120 stop_strong.n51 VSS 0.033109f
C2121 stop_strong.n52 VSS 0.049874f
C2122 stop_strong.n53 VSS 0.625244f
C2123 stop_strong.n54 VSS 0.558556f
C2124 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.936187f
C2125 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.087567f
C2126 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.039891f
C2127 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.097546f
C2128 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C2129 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C2130 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.115133f
C2131 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C2132 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.095888f
C2133 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.041221f
C2134 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C2135 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.108538f
C2136 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.081767f
C2137 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.090596f
C2138 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C2139 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.398296f
C2140 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.36504f
C2141 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C2142 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n7 VSS 0.753756f
C2143 a_3116_2192.t2 VSS 0.059028f
C2144 a_3116_2192.t5 VSS 0.059028f
C2145 a_3116_2192.t4 VSS 0.059028f
C2146 a_3116_2192.n0 VSS 0.139449f
C2147 a_3116_2192.t3 VSS 0.059028f
C2148 a_3116_2192.t1 VSS 0.059028f
C2149 a_3116_2192.n1 VSS 0.136068f
C2150 a_3116_2192.n2 VSS 1.11221f
C2151 a_3116_2192.n3 VSS 0.258102f
C2152 a_3116_2192.t0 VSS 0.059028f
C2153 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C2154 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.087824f
C2155 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.040008f
C2156 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C2157 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C2158 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.202807f
C2159 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.096169f
C2160 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.041341f
C2161 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C2162 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.082007f
C2163 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.090862f
C2164 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C2165 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C2166 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.107599f
C2167 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C2168 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C2169 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C2170 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C2171 saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
C2172 VDD.n0 VSS 0.097016f
C2173 VDD.t196 VSS 0.018573f
C2174 VDD.t236 VSS 0.018573f
C2175 VDD.n1 VSS 0.039357f
C2176 VDD.t271 VSS 0.070015f
C2177 VDD.n2 VSS 0.069693f
C2178 VDD.t19 VSS 0.070015f
C2179 VDD.n3 VSS 0.161184f
C2180 VDD.t198 VSS 0.018573f
C2181 VDD.t234 VSS 0.018573f
C2182 VDD.n4 VSS 0.039357f
C2183 VDD.n5 VSS 0.337883f
C2184 VDD.n6 VSS 0.114915f
C2185 VDD.n7 VSS 0.367811f
C2186 VDD.n8 VSS 0.139996f
C2187 VDD.t197 VSS 0.285918f
C2188 VDD.t233 VSS 0.180346f
C2189 VDD.t192 VSS 0.180346f
C2190 VDD.t18 VSS 0.236705f
C2191 VDD.n9 VSS 0.364397f
C2192 VDD.t235 VSS 0.280997f
C2193 VDD.t195 VSS 0.180346f
C2194 VDD.t265 VSS 0.180346f
C2195 VDD.t270 VSS 0.238754f
C2196 VDD.n10 VSS 0.042192f
C2197 VDD.n11 VSS 0.15063f
C2198 VDD.n12 VSS 0.148581f
C2199 VDD.n13 VSS 0.123157f
C2200 VDD.n14 VSS 0.139996f
C2201 VDD.n15 VSS 0.123157f
C2202 VDD.n16 VSS 0.010996f
C2203 VDD.n17 VSS 0.06159f
C2204 VDD.n18 VSS 0.161402f
C2205 VDD.n19 VSS 0.164495f
C2206 VDD.n20 VSS 0.08097f
C2207 VDD.n21 VSS 0.097153f
C2208 VDD.t277 VSS 0.018573f
C2209 VDD.t269 VSS 0.018573f
C2210 VDD.n22 VSS 0.039357f
C2211 VDD.t144 VSS 0.070015f
C2212 VDD.n23 VSS 0.06159f
C2213 VDD.n24 VSS 0.123157f
C2214 VDD.n25 VSS 0.069693f
C2215 VDD.t165 VSS 0.018573f
C2216 VDD.t71 VSS 0.018573f
C2217 VDD.n26 VSS 0.039357f
C2218 VDD.t218 VSS 0.070015f
C2219 VDD.n27 VSS 0.161402f
C2220 VDD.n28 VSS 0.164495f
C2221 VDD.n29 VSS 0.097153f
C2222 VDD.t97 VSS 0.018573f
C2223 VDD.t39 VSS 0.018573f
C2224 VDD.n30 VSS 0.039357f
C2225 VDD.t208 VSS 0.070015f
C2226 VDD.n31 VSS 0.06159f
C2227 VDD.n32 VSS 0.123157f
C2228 VDD.n33 VSS 0.069693f
C2229 VDD.t121 VSS 0.018573f
C2230 VDD.t41 VSS 0.018573f
C2231 VDD.n34 VSS 0.039357f
C2232 VDD.t163 VSS 0.070015f
C2233 VDD.n35 VSS 0.161402f
C2234 VDD.n36 VSS 0.164495f
C2235 VDD.n37 VSS 0.097153f
C2236 VDD.t172 VSS 0.018573f
C2237 VDD.t136 VSS 0.018573f
C2238 VDD.n38 VSS 0.039357f
C2239 VDD.t212 VSS 0.070015f
C2240 VDD.n39 VSS 0.06159f
C2241 VDD.n40 VSS 0.123157f
C2242 VDD.n41 VSS 0.069693f
C2243 VDD.t287 VSS 0.018573f
C2244 VDD.t91 VSS 0.018573f
C2245 VDD.n42 VSS 0.039357f
C2246 VDD.t127 VSS 0.070015f
C2247 VDD.n43 VSS 0.161402f
C2248 VDD.n44 VSS 0.164495f
C2249 VDD.n45 VSS 0.097153f
C2250 VDD.t27 VSS 0.018573f
C2251 VDD.t182 VSS 0.018573f
C2252 VDD.n46 VSS 0.039357f
C2253 VDD.t50 VSS 0.070015f
C2254 VDD.n47 VSS 0.06159f
C2255 VDD.n48 VSS 0.123157f
C2256 VDD.n49 VSS 0.069693f
C2257 VDD.t254 VSS 0.018573f
C2258 VDD.t223 VSS 0.018573f
C2259 VDD.n50 VSS 0.039357f
C2260 VDD.t267 VSS 0.070015f
C2261 VDD.n51 VSS 0.161402f
C2262 VDD.n52 VSS 0.164495f
C2263 VDD.n53 VSS 0.097153f
C2264 VDD.t59 VSS 0.018573f
C2265 VDD.t95 VSS 0.018573f
C2266 VDD.n54 VSS 0.039357f
C2267 VDD.t7 VSS 0.070015f
C2268 VDD.n55 VSS 0.06159f
C2269 VDD.n56 VSS 0.123157f
C2270 VDD.n57 VSS 0.069693f
C2271 VDD.t206 VSS 0.018573f
C2272 VDD.t230 VSS 0.018573f
C2273 VDD.n58 VSS 0.039357f
C2274 VDD.t47 VSS 0.070015f
C2275 VDD.n59 VSS 0.161402f
C2276 VDD.n60 VSS 0.164495f
C2277 VDD.n61 VSS 0.097153f
C2278 VDD.t103 VSS 0.018573f
C2279 VDD.t105 VSS 0.018573f
C2280 VDD.n62 VSS 0.039357f
C2281 VDD.t52 VSS 0.070015f
C2282 VDD.n63 VSS 0.06159f
C2283 VDD.n64 VSS 0.123157f
C2284 VDD.n65 VSS 0.069693f
C2285 VDD.t140 VSS 0.018573f
C2286 VDD.t63 VSS 0.018573f
C2287 VDD.n66 VSS 0.039357f
C2288 VDD.t216 VSS 0.070015f
C2289 VDD.n67 VSS 0.161402f
C2290 VDD.n68 VSS 0.164495f
C2291 VDD.n69 VSS 0.097153f
C2292 VDD.t61 VSS 0.018573f
C2293 VDD.t5 VSS 0.018573f
C2294 VDD.n70 VSS 0.039357f
C2295 VDD.t301 VSS 0.070015f
C2296 VDD.n71 VSS 0.06159f
C2297 VDD.n72 VSS 0.123157f
C2298 VDD.n73 VSS 0.069693f
C2299 VDD.t260 VSS 0.018573f
C2300 VDD.t293 VSS 0.018573f
C2301 VDD.n74 VSS 0.039357f
C2302 VDD.t295 VSS 0.070015f
C2303 VDD.n75 VSS 0.161402f
C2304 VDD.n76 VSS 0.164495f
C2305 VDD.n77 VSS 0.09525f
C2306 VDD.t154 VSS 0.069612f
C2307 VDD.t37 VSS 0.069612f
C2308 VDD.t138 VSS 0.069612f
C2309 VDD.t279 VSS 0.070299f
C2310 VDD.n78 VSS 0.259059f
C2311 VDD.n79 VSS 0.137385f
C2312 VDD.n80 VSS 0.128449f
C2313 VDD.n81 VSS 0.09525f
C2314 VDD.t107 VSS 0.069612f
C2315 VDD.t291 VSS 0.069612f
C2316 VDD.t123 VSS 0.069612f
C2317 VDD.t109 VSS 0.070299f
C2318 VDD.n82 VSS 0.259059f
C2319 VDD.n83 VSS 0.137385f
C2320 VDD.n84 VSS 0.128449f
C2321 VDD.n85 VSS 0.09525f
C2322 VDD.t174 VSS 0.069612f
C2323 VDD.t210 VSS 0.069612f
C2324 VDD.t31 VSS 0.069612f
C2325 VDD.t214 VSS 0.070299f
C2326 VDD.n86 VSS 0.259059f
C2327 VDD.n87 VSS 0.137385f
C2328 VDD.n88 VSS 0.128449f
C2329 VDD.n89 VSS 0.09525f
C2330 VDD.t156 VSS 0.069612f
C2331 VDD.t134 VSS 0.069612f
C2332 VDD.t315 VSS 0.069612f
C2333 VDD.t23 VSS 0.070299f
C2334 VDD.n90 VSS 0.259059f
C2335 VDD.n91 VSS 0.137385f
C2336 VDD.n92 VSS 0.128449f
C2337 VDD.n93 VSS 0.09525f
C2338 VDD.t93 VSS 0.069612f
C2339 VDD.t303 VSS 0.069612f
C2340 VDD.t119 VSS 0.069612f
C2341 VDD.t21 VSS 0.070299f
C2342 VDD.n94 VSS 0.259059f
C2343 VDD.n95 VSS 0.137385f
C2344 VDD.n96 VSS 0.128449f
C2345 VDD.n97 VSS 0.09525f
C2346 VDD.t309 VSS 0.069612f
C2347 VDD.t43 VSS 0.069612f
C2348 VDD.t148 VSS 0.069612f
C2349 VDD.t311 VSS 0.070299f
C2350 VDD.n98 VSS 0.259059f
C2351 VDD.n99 VSS 0.137385f
C2352 VDD.n100 VSS 0.128449f
C2353 VDD.n101 VSS 0.09525f
C2354 VDD.t9 VSS 0.069612f
C2355 VDD.t180 VSS 0.069612f
C2356 VDD.t150 VSS 0.069612f
C2357 VDD.t262 VSS 0.070299f
C2358 VDD.n102 VSS 0.259059f
C2359 VDD.n103 VSS 0.137385f
C2360 VDD.n104 VSS 0.128449f
C2361 VDD.n105 VSS 0.09525f
C2362 VDD.t125 VSS 0.069612f
C2363 VDD.t232 VSS 0.069612f
C2364 VDD.t194 VSS 0.069612f
C2365 VDD.t152 VSS 0.070299f
C2366 VDD.n106 VSS 0.259059f
C2367 VDD.n107 VSS 0.137385f
C2368 VDD.n108 VSS 0.128449f
C2369 VDD.n109 VSS 0.435069f
C2370 VDD.n110 VSS 0.391663f
C2371 VDD.t151 VSS 0.301961f
C2372 VDD.t193 VSS 0.333897f
C2373 VDD.n111 VSS 0.249855f
C2374 VDD.n112 VSS 0.319044f
C2375 VDD.t124 VSS 0.298176f
C2376 VDD.t231 VSS 0.349797f
C2377 VDD.n113 VSS 0.684675f
C2378 VDD.n114 VSS 0.065409f
C2379 VDD.n115 VSS 0.658688f
C2380 VDD.n116 VSS 0.364449f
C2381 VDD.n117 VSS 0.149291f
C2382 VDD.n118 VSS 0.435069f
C2383 VDD.n119 VSS 0.391663f
C2384 VDD.t261 VSS 0.301961f
C2385 VDD.t149 VSS 0.333897f
C2386 VDD.n120 VSS 0.249855f
C2387 VDD.n121 VSS 0.319044f
C2388 VDD.t8 VSS 0.298176f
C2389 VDD.t179 VSS 0.349797f
C2390 VDD.n122 VSS 0.684675f
C2391 VDD.n123 VSS 0.065409f
C2392 VDD.n124 VSS 0.432347f
C2393 VDD.n125 VSS 0.283834f
C2394 VDD.n126 VSS 0.084847f
C2395 VDD.n127 VSS 0.149291f
C2396 VDD.n128 VSS 0.435069f
C2397 VDD.n129 VSS 0.391663f
C2398 VDD.t310 VSS 0.301961f
C2399 VDD.t147 VSS 0.333897f
C2400 VDD.n130 VSS 0.249855f
C2401 VDD.n131 VSS 0.319044f
C2402 VDD.t308 VSS 0.298176f
C2403 VDD.t42 VSS 0.349797f
C2404 VDD.n132 VSS 0.684675f
C2405 VDD.n133 VSS 0.065409f
C2406 VDD.n134 VSS 0.432347f
C2407 VDD.n135 VSS 0.283834f
C2408 VDD.n136 VSS 0.084847f
C2409 VDD.n137 VSS 0.149291f
C2410 VDD.n138 VSS 0.435069f
C2411 VDD.n139 VSS 0.391663f
C2412 VDD.t20 VSS 0.301961f
C2413 VDD.t118 VSS 0.333897f
C2414 VDD.n140 VSS 0.249855f
C2415 VDD.n141 VSS 0.319044f
C2416 VDD.t92 VSS 0.298176f
C2417 VDD.t302 VSS 0.349797f
C2418 VDD.n142 VSS 0.684675f
C2419 VDD.n143 VSS 0.065409f
C2420 VDD.n144 VSS 0.432347f
C2421 VDD.n145 VSS 0.283834f
C2422 VDD.n146 VSS 0.084847f
C2423 VDD.n147 VSS 0.149291f
C2424 VDD.n148 VSS 0.435069f
C2425 VDD.n149 VSS 0.391663f
C2426 VDD.t22 VSS 0.301961f
C2427 VDD.t314 VSS 0.333897f
C2428 VDD.n150 VSS 0.249855f
C2429 VDD.n151 VSS 0.319044f
C2430 VDD.t155 VSS 0.298176f
C2431 VDD.t133 VSS 0.349797f
C2432 VDD.n152 VSS 0.684675f
C2433 VDD.n153 VSS 0.065409f
C2434 VDD.n154 VSS 0.432347f
C2435 VDD.n155 VSS 0.283834f
C2436 VDD.n156 VSS 0.084847f
C2437 VDD.n157 VSS 0.149291f
C2438 VDD.n158 VSS 0.435069f
C2439 VDD.n159 VSS 0.391663f
C2440 VDD.t213 VSS 0.301961f
C2441 VDD.t30 VSS 0.333897f
C2442 VDD.n160 VSS 0.249855f
C2443 VDD.n161 VSS 0.319044f
C2444 VDD.t173 VSS 0.298176f
C2445 VDD.t209 VSS 0.349797f
C2446 VDD.n162 VSS 0.684675f
C2447 VDD.n163 VSS 0.065409f
C2448 VDD.n164 VSS 0.432347f
C2449 VDD.n165 VSS 0.283834f
C2450 VDD.n166 VSS 0.084847f
C2451 VDD.n167 VSS 0.149291f
C2452 VDD.n168 VSS 0.435069f
C2453 VDD.n169 VSS 0.391663f
C2454 VDD.t108 VSS 0.301961f
C2455 VDD.t122 VSS 0.333897f
C2456 VDD.n170 VSS 0.249855f
C2457 VDD.n171 VSS 0.319044f
C2458 VDD.t106 VSS 0.298176f
C2459 VDD.t290 VSS 0.349797f
C2460 VDD.n172 VSS 0.684675f
C2461 VDD.n173 VSS 0.065409f
C2462 VDD.n174 VSS 0.432347f
C2463 VDD.n175 VSS 0.283834f
C2464 VDD.n176 VSS 0.084847f
C2465 VDD.n177 VSS 0.149291f
C2466 VDD.n178 VSS 0.435069f
C2467 VDD.n179 VSS 0.391663f
C2468 VDD.t278 VSS 0.301961f
C2469 VDD.t137 VSS 0.333897f
C2470 VDD.n180 VSS 0.249855f
C2471 VDD.n181 VSS 0.319044f
C2472 VDD.t153 VSS 0.298176f
C2473 VDD.t36 VSS 0.349797f
C2474 VDD.n182 VSS 0.684675f
C2475 VDD.n183 VSS 0.065409f
C2476 VDD.n184 VSS 0.432347f
C2477 VDD.n185 VSS 0.283834f
C2478 VDD.n186 VSS 0.084847f
C2479 VDD.n187 VSS 0.149291f
C2480 VDD.n188 VSS 0.109134f
C2481 VDD.t281 VSS 0.018573f
C2482 VDD.t67 VSS 0.018573f
C2483 VDD.n189 VSS 0.0397f
C2484 VDD.t275 VSS 0.018573f
C2485 VDD.t202 VSS 0.018573f
C2486 VDD.n190 VSS 0.0397f
C2487 VDD.t244 VSS 0.018573f
C2488 VDD.t240 VSS 0.018573f
C2489 VDD.n191 VSS 0.0397f
C2490 VDD.n192 VSS 0.160193f
C2491 VDD.n193 VSS 0.098311f
C2492 VDD.n194 VSS 0.109134f
C2493 VDD.t252 VSS 0.018573f
C2494 VDD.t250 VSS 0.018573f
C2495 VDD.n195 VSS 0.0397f
C2496 VDD.t248 VSS 0.018573f
C2497 VDD.t246 VSS 0.018573f
C2498 VDD.n196 VSS 0.0397f
C2499 VDD.t75 VSS 0.018573f
C2500 VDD.t81 VSS 0.018573f
C2501 VDD.n197 VSS 0.0397f
C2502 VDD.n198 VSS 0.160193f
C2503 VDD.n199 VSS 0.098311f
C2504 VDD.n200 VSS 0.109134f
C2505 VDD.t3 VSS 0.018573f
C2506 VDD.t15 VSS 0.018573f
C2507 VDD.n201 VSS 0.0397f
C2508 VDD.t17 VSS 0.018573f
C2509 VDD.t1 VSS 0.018573f
C2510 VDD.n202 VSS 0.0397f
C2511 VDD.t191 VSS 0.018573f
C2512 VDD.t87 VSS 0.018573f
C2513 VDD.n203 VSS 0.0397f
C2514 VDD.n204 VSS 0.160193f
C2515 VDD.n205 VSS 0.098311f
C2516 VDD.n206 VSS 0.109134f
C2517 VDD.t319 VSS 0.018573f
C2518 VDD.t83 VSS 0.018573f
C2519 VDD.n207 VSS 0.0397f
C2520 VDD.t317 VSS 0.018573f
C2521 VDD.t273 VSS 0.018573f
C2522 VDD.n208 VSS 0.0397f
C2523 VDD.t220 VSS 0.018573f
C2524 VDD.t200 VSS 0.018573f
C2525 VDD.n209 VSS 0.0397f
C2526 VDD.n210 VSS 0.160193f
C2527 VDD.n211 VSS 0.098311f
C2528 VDD.n212 VSS 0.109134f
C2529 VDD.t176 VSS 0.018573f
C2530 VDD.t65 VSS 0.018573f
C2531 VDD.n213 VSS 0.0397f
C2532 VDD.t55 VSS 0.018573f
C2533 VDD.t25 VSS 0.018573f
C2534 VDD.n214 VSS 0.0397f
C2535 VDD.t204 VSS 0.018573f
C2536 VDD.t264 VSS 0.018573f
C2537 VDD.n215 VSS 0.0397f
C2538 VDD.n216 VSS 0.160193f
C2539 VDD.n217 VSS 0.098311f
C2540 VDD.n218 VSS 0.109134f
C2541 VDD.t285 VSS 0.018573f
C2542 VDD.t313 VSS 0.018573f
C2543 VDD.n219 VSS 0.0397f
C2544 VDD.t111 VSS 0.018573f
C2545 VDD.t132 VSS 0.018573f
C2546 VDD.n220 VSS 0.0397f
C2547 VDD.t228 VSS 0.018573f
C2548 VDD.t283 VSS 0.018573f
C2549 VDD.n221 VSS 0.0397f
C2550 VDD.n222 VSS 0.160193f
C2551 VDD.n223 VSS 0.098311f
C2552 VDD.n224 VSS 0.109134f
C2553 VDD.t161 VSS 0.018573f
C2554 VDD.t29 VSS 0.018573f
C2555 VDD.n225 VSS 0.0397f
C2556 VDD.t57 VSS 0.018573f
C2557 VDD.t99 VSS 0.018573f
C2558 VDD.n226 VSS 0.0397f
C2559 VDD.t258 VSS 0.018573f
C2560 VDD.t307 VSS 0.018573f
C2561 VDD.n227 VSS 0.0397f
C2562 VDD.n228 VSS 0.160193f
C2563 VDD.n229 VSS 0.098311f
C2564 VDD.n230 VSS 0.109134f
C2565 VDD.t35 VSS 0.018573f
C2566 VDD.t115 VSS 0.018573f
C2567 VDD.n231 VSS 0.0397f
C2568 VDD.t305 VSS 0.018573f
C2569 VDD.t289 VSS 0.018573f
C2570 VDD.n232 VSS 0.0397f
C2571 VDD.t187 VSS 0.018573f
C2572 VDD.t73 VSS 0.018573f
C2573 VDD.n233 VSS 0.0397f
C2574 VDD.n234 VSS 0.160193f
C2575 VDD.n235 VSS 0.098311f
C2576 VDD.n236 VSS 0.109134f
C2577 VDD.t117 VSS 0.018573f
C2578 VDD.t89 VSS 0.018573f
C2579 VDD.n237 VSS 0.0397f
C2580 VDD.t33 VSS 0.018573f
C2581 VDD.t256 VSS 0.018573f
C2582 VDD.n238 VSS 0.0397f
C2583 VDD.t12 VSS 0.018573f
C2584 VDD.t130 VSS 0.018573f
C2585 VDD.n239 VSS 0.0397f
C2586 VDD.n240 VSS 0.160193f
C2587 VDD.n241 VSS 0.098311f
C2588 VDD.t167 VSS 0.018573f
C2589 VDD.t69 VSS 0.018573f
C2590 VDD.n242 VSS 0.0397f
C2591 VDD.n243 VSS 0.230443f
C2592 VDD.n244 VSS 0.118188f
C2593 VDD.n245 VSS 0.12677f
C2594 VDD.n246 VSS 0.442174f
C2595 VDD.n247 VSS 0.321258f
C2596 VDD.t166 VSS 0.281899f
C2597 VDD.t68 VSS 0.191618f
C2598 VDD.t11 VSS 0.191618f
C2599 VDD.t129 VSS 0.254765f
C2600 VDD.n248 VSS 0.163311f
C2601 VDD.t88 VSS 0.295731f
C2602 VDD.t116 VSS 0.191618f
C2603 VDD.t255 VSS 0.191618f
C2604 VDD.t32 VSS 0.25041f
C2605 VDD.n249 VSS 0.158956f
C2606 VDD.n250 VSS 0.108723f
C2607 VDD.n251 VSS 0.108723f
C2608 VDD.n252 VSS 0.131726f
C2609 VDD.n253 VSS 0.038938f
C2610 VDD.n254 VSS 0.160193f
C2611 VDD.n255 VSS 0.16009f
C2612 VDD.n256 VSS 0.073617f
C2613 VDD.t299 VSS 0.018573f
C2614 VDD.t170 VSS 0.018573f
C2615 VDD.n257 VSS 0.0397f
C2616 VDD.n258 VSS 0.16009f
C2617 VDD.n259 VSS 0.182645f
C2618 VDD.n260 VSS 0.10939f
C2619 VDD.n261 VSS 0.12677f
C2620 VDD.n262 VSS 0.442174f
C2621 VDD.n263 VSS 0.321258f
C2622 VDD.t298 VSS 0.281899f
C2623 VDD.t169 VSS 0.191618f
C2624 VDD.t186 VSS 0.191618f
C2625 VDD.t72 VSS 0.254765f
C2626 VDD.n264 VSS 0.163311f
C2627 VDD.t114 VSS 0.295731f
C2628 VDD.t34 VSS 0.191618f
C2629 VDD.t288 VSS 0.191618f
C2630 VDD.t304 VSS 0.25041f
C2631 VDD.n265 VSS 0.158956f
C2632 VDD.n266 VSS 0.108723f
C2633 VDD.n267 VSS 0.108723f
C2634 VDD.n268 VSS 0.131726f
C2635 VDD.n269 VSS 0.038938f
C2636 VDD.n270 VSS 0.160193f
C2637 VDD.n271 VSS 0.16009f
C2638 VDD.n272 VSS 0.073617f
C2639 VDD.t146 VSS 0.018573f
C2640 VDD.t101 VSS 0.018573f
C2641 VDD.n273 VSS 0.0397f
C2642 VDD.n274 VSS 0.16009f
C2643 VDD.n275 VSS 0.182645f
C2644 VDD.n276 VSS 0.10939f
C2645 VDD.n277 VSS 0.12677f
C2646 VDD.n278 VSS 0.442174f
C2647 VDD.n279 VSS 0.321258f
C2648 VDD.t145 VSS 0.281899f
C2649 VDD.t100 VSS 0.191618f
C2650 VDD.t257 VSS 0.191618f
C2651 VDD.t306 VSS 0.254765f
C2652 VDD.n280 VSS 0.163311f
C2653 VDD.t28 VSS 0.295731f
C2654 VDD.t160 VSS 0.191618f
C2655 VDD.t98 VSS 0.191618f
C2656 VDD.t56 VSS 0.25041f
C2657 VDD.n281 VSS 0.158956f
C2658 VDD.n282 VSS 0.108723f
C2659 VDD.n283 VSS 0.108723f
C2660 VDD.n284 VSS 0.131726f
C2661 VDD.n285 VSS 0.038938f
C2662 VDD.n286 VSS 0.160193f
C2663 VDD.n287 VSS 0.16009f
C2664 VDD.n288 VSS 0.073617f
C2665 VDD.t226 VSS 0.018573f
C2666 VDD.t297 VSS 0.018573f
C2667 VDD.n289 VSS 0.0397f
C2668 VDD.n290 VSS 0.16009f
C2669 VDD.n291 VSS 0.182645f
C2670 VDD.n292 VSS 0.10939f
C2671 VDD.n293 VSS 0.12677f
C2672 VDD.n294 VSS 0.442174f
C2673 VDD.n295 VSS 0.321258f
C2674 VDD.t225 VSS 0.281899f
C2675 VDD.t296 VSS 0.191618f
C2676 VDD.t227 VSS 0.191618f
C2677 VDD.t282 VSS 0.254765f
C2678 VDD.n296 VSS 0.163311f
C2679 VDD.t312 VSS 0.295731f
C2680 VDD.t284 VSS 0.191618f
C2681 VDD.t131 VSS 0.191618f
C2682 VDD.t110 VSS 0.25041f
C2683 VDD.n297 VSS 0.158956f
C2684 VDD.n298 VSS 0.108723f
C2685 VDD.n299 VSS 0.108723f
C2686 VDD.n300 VSS 0.131726f
C2687 VDD.n301 VSS 0.038938f
C2688 VDD.n302 VSS 0.160193f
C2689 VDD.n303 VSS 0.16009f
C2690 VDD.n304 VSS 0.073617f
C2691 VDD.t185 VSS 0.018573f
C2692 VDD.t142 VSS 0.018573f
C2693 VDD.n305 VSS 0.0397f
C2694 VDD.n306 VSS 0.16009f
C2695 VDD.n307 VSS 0.182645f
C2696 VDD.n308 VSS 0.10939f
C2697 VDD.n309 VSS 0.12677f
C2698 VDD.n310 VSS 0.442174f
C2699 VDD.n311 VSS 0.321258f
C2700 VDD.t184 VSS 0.281899f
C2701 VDD.t141 VSS 0.191618f
C2702 VDD.t203 VSS 0.191618f
C2703 VDD.t263 VSS 0.254765f
C2704 VDD.n312 VSS 0.163311f
C2705 VDD.t64 VSS 0.295731f
C2706 VDD.t175 VSS 0.191618f
C2707 VDD.t24 VSS 0.191618f
C2708 VDD.t54 VSS 0.25041f
C2709 VDD.n313 VSS 0.158956f
C2710 VDD.n314 VSS 0.108723f
C2711 VDD.n315 VSS 0.108723f
C2712 VDD.n316 VSS 0.131726f
C2713 VDD.n317 VSS 0.038938f
C2714 VDD.n318 VSS 0.160193f
C2715 VDD.n319 VSS 0.16009f
C2716 VDD.n320 VSS 0.073617f
C2717 VDD.t113 VSS 0.018573f
C2718 VDD.t189 VSS 0.018573f
C2719 VDD.n321 VSS 0.0397f
C2720 VDD.n322 VSS 0.16009f
C2721 VDD.n323 VSS 0.182645f
C2722 VDD.n324 VSS 0.10939f
C2723 VDD.n325 VSS 0.12677f
C2724 VDD.n326 VSS 0.442174f
C2725 VDD.n327 VSS 0.321258f
C2726 VDD.t112 VSS 0.281899f
C2727 VDD.t188 VSS 0.191618f
C2728 VDD.t219 VSS 0.191618f
C2729 VDD.t199 VSS 0.254765f
C2730 VDD.n328 VSS 0.163311f
C2731 VDD.t82 VSS 0.295731f
C2732 VDD.t318 VSS 0.191618f
C2733 VDD.t272 VSS 0.191618f
C2734 VDD.t316 VSS 0.25041f
C2735 VDD.n329 VSS 0.158956f
C2736 VDD.n330 VSS 0.108723f
C2737 VDD.n331 VSS 0.108723f
C2738 VDD.n332 VSS 0.131726f
C2739 VDD.n333 VSS 0.038938f
C2740 VDD.n334 VSS 0.160193f
C2741 VDD.n335 VSS 0.16009f
C2742 VDD.n336 VSS 0.073617f
C2743 VDD.t178 VSS 0.018573f
C2744 VDD.t85 VSS 0.018573f
C2745 VDD.n337 VSS 0.0397f
C2746 VDD.n338 VSS 0.16009f
C2747 VDD.n339 VSS 0.182645f
C2748 VDD.n340 VSS 0.10939f
C2749 VDD.n341 VSS 0.12677f
C2750 VDD.n342 VSS 0.442174f
C2751 VDD.n343 VSS 0.321258f
C2752 VDD.t177 VSS 0.281899f
C2753 VDD.t84 VSS 0.191618f
C2754 VDD.t190 VSS 0.191618f
C2755 VDD.t86 VSS 0.254765f
C2756 VDD.n344 VSS 0.163311f
C2757 VDD.t14 VSS 0.295731f
C2758 VDD.t2 VSS 0.191618f
C2759 VDD.t0 VSS 0.191618f
C2760 VDD.t16 VSS 0.25041f
C2761 VDD.n345 VSS 0.158956f
C2762 VDD.n346 VSS 0.108723f
C2763 VDD.n347 VSS 0.108723f
C2764 VDD.n348 VSS 0.131726f
C2765 VDD.n349 VSS 0.038938f
C2766 VDD.n350 VSS 0.160193f
C2767 VDD.n351 VSS 0.16009f
C2768 VDD.n352 VSS 0.073617f
C2769 VDD.t77 VSS 0.018573f
C2770 VDD.t79 VSS 0.018573f
C2771 VDD.n353 VSS 0.0397f
C2772 VDD.n354 VSS 0.16009f
C2773 VDD.n355 VSS 0.182645f
C2774 VDD.n356 VSS 0.10939f
C2775 VDD.n357 VSS 0.12677f
C2776 VDD.n358 VSS 0.442174f
C2777 VDD.n359 VSS 0.321258f
C2778 VDD.t76 VSS 0.281899f
C2779 VDD.t78 VSS 0.191618f
C2780 VDD.t74 VSS 0.191618f
C2781 VDD.t80 VSS 0.254765f
C2782 VDD.n360 VSS 0.163311f
C2783 VDD.t249 VSS 0.295731f
C2784 VDD.t251 VSS 0.191618f
C2785 VDD.t245 VSS 0.191618f
C2786 VDD.t247 VSS 0.25041f
C2787 VDD.n361 VSS 0.158956f
C2788 VDD.n362 VSS 0.108723f
C2789 VDD.n363 VSS 0.108723f
C2790 VDD.n364 VSS 0.131726f
C2791 VDD.n365 VSS 0.038938f
C2792 VDD.n366 VSS 0.160193f
C2793 VDD.n367 VSS 0.16009f
C2794 VDD.n368 VSS 0.073617f
C2795 VDD.t242 VSS 0.018573f
C2796 VDD.t238 VSS 0.018573f
C2797 VDD.n369 VSS 0.0397f
C2798 VDD.n370 VSS 0.16009f
C2799 VDD.n371 VSS 0.182645f
C2800 VDD.n372 VSS 0.10939f
C2801 VDD.n373 VSS 0.12677f
C2802 VDD.n374 VSS 0.442174f
C2803 VDD.n375 VSS 0.321258f
C2804 VDD.t241 VSS 0.281899f
C2805 VDD.t237 VSS 0.191618f
C2806 VDD.t243 VSS 0.191618f
C2807 VDD.t239 VSS 0.254765f
C2808 VDD.n376 VSS 0.163311f
C2809 VDD.t66 VSS 0.295731f
C2810 VDD.t280 VSS 0.191618f
C2811 VDD.t201 VSS 0.191618f
C2812 VDD.t274 VSS 0.25041f
C2813 VDD.n377 VSS 0.158956f
C2814 VDD.n378 VSS 0.108723f
C2815 VDD.n379 VSS 0.108723f
C2816 VDD.n380 VSS 0.131726f
C2817 VDD.n381 VSS 0.038938f
C2818 VDD.n382 VSS 0.160193f
C2819 VDD.n383 VSS 0.16009f
C2820 VDD.n384 VSS 0.073617f
C2821 VDD.n385 VSS 1.02788f
C2822 VDD.n386 VSS 0.08097f
C2823 VDD.n387 VSS 0.139996f
C2824 VDD.n388 VSS 0.367811f
C2825 VDD.t60 VSS 0.285918f
C2826 VDD.t4 VSS 0.180346f
C2827 VDD.t44 VSS 0.180346f
C2828 VDD.t300 VSS 0.236705f
C2829 VDD.n389 VSS 0.148581f
C2830 VDD.n390 VSS 0.042192f
C2831 VDD.n391 VSS 0.15063f
C2832 VDD.t294 VSS 0.238754f
C2833 VDD.t45 VSS 0.180346f
C2834 VDD.t259 VSS 0.180346f
C2835 VDD.t292 VSS 0.280997f
C2836 VDD.n392 VSS 0.364397f
C2837 VDD.n393 VSS 0.097016f
C2838 VDD.n394 VSS 0.139996f
C2839 VDD.n395 VSS 0.123157f
C2840 VDD.n396 VSS 0.010996f
C2841 VDD.n397 VSS 0.161184f
C2842 VDD.n398 VSS 0.165148f
C2843 VDD.n399 VSS 0.131052f
C2844 VDD.n400 VSS 0.08097f
C2845 VDD.n401 VSS 0.139996f
C2846 VDD.n402 VSS 0.367811f
C2847 VDD.t102 VSS 0.285918f
C2848 VDD.t104 VSS 0.180346f
C2849 VDD.t53 VSS 0.180346f
C2850 VDD.t51 VSS 0.236705f
C2851 VDD.n403 VSS 0.148581f
C2852 VDD.n404 VSS 0.042192f
C2853 VDD.n405 VSS 0.15063f
C2854 VDD.t215 VSS 0.238754f
C2855 VDD.t48 VSS 0.180346f
C2856 VDD.t139 VSS 0.180346f
C2857 VDD.t62 VSS 0.280997f
C2858 VDD.n406 VSS 0.364397f
C2859 VDD.n407 VSS 0.097016f
C2860 VDD.n408 VSS 0.139996f
C2861 VDD.n409 VSS 0.123157f
C2862 VDD.n410 VSS 0.010996f
C2863 VDD.n411 VSS 0.161184f
C2864 VDD.n412 VSS 0.165148f
C2865 VDD.n413 VSS 0.131052f
C2866 VDD.n414 VSS 0.08097f
C2867 VDD.n415 VSS 0.139996f
C2868 VDD.n416 VSS 0.367811f
C2869 VDD.t58 VSS 0.285918f
C2870 VDD.t94 VSS 0.180346f
C2871 VDD.t159 VSS 0.180346f
C2872 VDD.t6 VSS 0.236705f
C2873 VDD.n417 VSS 0.148581f
C2874 VDD.n418 VSS 0.042192f
C2875 VDD.n419 VSS 0.15063f
C2876 VDD.t46 VSS 0.238754f
C2877 VDD.t224 VSS 0.180346f
C2878 VDD.t205 VSS 0.180346f
C2879 VDD.t229 VSS 0.280997f
C2880 VDD.n420 VSS 0.364397f
C2881 VDD.n421 VSS 0.097016f
C2882 VDD.n422 VSS 0.139996f
C2883 VDD.n423 VSS 0.123157f
C2884 VDD.n424 VSS 0.010996f
C2885 VDD.n425 VSS 0.161184f
C2886 VDD.n426 VSS 0.165148f
C2887 VDD.n427 VSS 0.131052f
C2888 VDD.n428 VSS 0.08097f
C2889 VDD.n429 VSS 0.139996f
C2890 VDD.n430 VSS 0.367811f
C2891 VDD.t26 VSS 0.285918f
C2892 VDD.t181 VSS 0.180346f
C2893 VDD.t168 VSS 0.180346f
C2894 VDD.t49 VSS 0.236705f
C2895 VDD.n431 VSS 0.148581f
C2896 VDD.n432 VSS 0.042192f
C2897 VDD.n433 VSS 0.15063f
C2898 VDD.t266 VSS 0.238754f
C2899 VDD.t158 VSS 0.180346f
C2900 VDD.t253 VSS 0.180346f
C2901 VDD.t222 VSS 0.280997f
C2902 VDD.n434 VSS 0.364397f
C2903 VDD.n435 VSS 0.097016f
C2904 VDD.n436 VSS 0.139996f
C2905 VDD.n437 VSS 0.123157f
C2906 VDD.n438 VSS 0.010996f
C2907 VDD.n439 VSS 0.161184f
C2908 VDD.n440 VSS 0.165148f
C2909 VDD.n441 VSS 0.131052f
C2910 VDD.n442 VSS 0.08097f
C2911 VDD.n443 VSS 0.139996f
C2912 VDD.n444 VSS 0.367811f
C2913 VDD.t171 VSS 0.285918f
C2914 VDD.t135 VSS 0.180346f
C2915 VDD.t128 VSS 0.180346f
C2916 VDD.t211 VSS 0.236705f
C2917 VDD.n445 VSS 0.148581f
C2918 VDD.n446 VSS 0.042192f
C2919 VDD.n447 VSS 0.15063f
C2920 VDD.t126 VSS 0.238754f
C2921 VDD.t13 VSS 0.180346f
C2922 VDD.t286 VSS 0.180346f
C2923 VDD.t90 VSS 0.280997f
C2924 VDD.n448 VSS 0.364397f
C2925 VDD.n449 VSS 0.097016f
C2926 VDD.n450 VSS 0.139996f
C2927 VDD.n451 VSS 0.123157f
C2928 VDD.n452 VSS 0.010996f
C2929 VDD.n453 VSS 0.161184f
C2930 VDD.n454 VSS 0.165148f
C2931 VDD.n455 VSS 0.131052f
C2932 VDD.n456 VSS 0.08097f
C2933 VDD.n457 VSS 0.139996f
C2934 VDD.n458 VSS 0.367811f
C2935 VDD.t96 VSS 0.285918f
C2936 VDD.t38 VSS 0.180346f
C2937 VDD.t221 VSS 0.180346f
C2938 VDD.t207 VSS 0.236705f
C2939 VDD.n459 VSS 0.148581f
C2940 VDD.n460 VSS 0.042192f
C2941 VDD.n461 VSS 0.15063f
C2942 VDD.t162 VSS 0.238754f
C2943 VDD.t157 VSS 0.180346f
C2944 VDD.t120 VSS 0.180346f
C2945 VDD.t40 VSS 0.280997f
C2946 VDD.n462 VSS 0.364397f
C2947 VDD.n463 VSS 0.097016f
C2948 VDD.n464 VSS 0.139996f
C2949 VDD.n465 VSS 0.123157f
C2950 VDD.n466 VSS 0.010996f
C2951 VDD.n467 VSS 0.161184f
C2952 VDD.n468 VSS 0.165148f
C2953 VDD.n469 VSS 0.131052f
C2954 VDD.n470 VSS 0.08097f
C2955 VDD.n471 VSS 0.139996f
C2956 VDD.n472 VSS 0.367811f
C2957 VDD.t276 VSS 0.285918f
C2958 VDD.t268 VSS 0.180346f
C2959 VDD.t10 VSS 0.180346f
C2960 VDD.t143 VSS 0.236705f
C2961 VDD.n473 VSS 0.148581f
C2962 VDD.n474 VSS 0.042192f
C2963 VDD.n475 VSS 0.15063f
C2964 VDD.t217 VSS 0.238754f
C2965 VDD.t183 VSS 0.180346f
C2966 VDD.t164 VSS 0.180346f
C2967 VDD.t70 VSS 0.280997f
C2968 VDD.n476 VSS 0.364397f
C2969 VDD.n477 VSS 0.097016f
C2970 VDD.n478 VSS 0.139996f
C2971 VDD.n479 VSS 0.123157f
C2972 VDD.n480 VSS 0.010996f
C2973 VDD.n481 VSS 0.161184f
C2974 VDD.n482 VSS 0.165148f
C2975 VDD.n483 VSS 0.131052f
C2976 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C2977 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.087824f
C2978 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.040008f
C2979 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C2980 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C2981 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.202807f
C2982 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.096169f
C2983 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.041341f
C2984 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C2985 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.082007f
C2986 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.090862f
C2987 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C2988 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C2989 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.107599f
C2990 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C2991 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C2992 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C2993 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C2994 saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
.ends

