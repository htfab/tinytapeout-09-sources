`ifndef LOGO_NAME
`define LOGO_NAME logo
`endif
`ifndef LOGO_INSTANCE
`define LOGO_INSTANCE um_logo
`endif

(* blackbox *)
module `LOGO_NAME ();
endmodule
