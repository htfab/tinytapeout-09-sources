magic
tech sky130A
magscale 1 2
timestamp 1729594661
<< error_p >>
rect -31 272 31 278
rect -31 238 -19 272
rect -31 232 31 238
rect -31 -238 31 -232
rect -31 -272 -19 -238
rect -31 -278 31 -272
<< pwell >>
rect -231 -410 231 410
<< nmoslvt >>
rect -35 -200 35 200
<< ndiff >>
rect -93 188 -35 200
rect -93 -188 -81 188
rect -47 -188 -35 188
rect -93 -200 -35 -188
rect 35 188 93 200
rect 35 -188 47 188
rect 81 -188 93 188
rect 35 -200 93 -188
<< ndiffc >>
rect -81 -188 -47 188
rect 47 -188 81 188
<< psubdiff >>
rect -195 340 -99 374
rect 99 340 195 374
rect -195 278 -161 340
rect 161 278 195 340
rect -195 -340 -161 -278
rect 161 -340 195 -278
rect -195 -374 -99 -340
rect 99 -374 195 -340
<< psubdiffcont >>
rect -99 340 99 374
rect -195 -278 -161 278
rect 161 -278 195 278
rect -99 -374 99 -340
<< poly >>
rect -35 272 35 288
rect -35 238 -19 272
rect 19 238 35 272
rect -35 200 35 238
rect -35 -238 35 -200
rect -35 -272 -19 -238
rect 19 -272 35 -238
rect -35 -288 35 -272
<< polycont >>
rect -19 238 19 272
rect -19 -272 19 -238
<< locali >>
rect -195 340 -99 374
rect 99 340 195 374
rect -195 278 -161 340
rect 161 278 195 340
rect -35 238 -19 272
rect 19 238 35 272
rect -81 188 -47 204
rect -81 -204 -47 -188
rect 47 188 81 204
rect 47 -204 81 -188
rect -35 -272 -19 -238
rect 19 -272 35 -238
rect -195 -340 -161 -278
rect 161 -340 195 -278
rect -195 -374 -99 -340
rect 99 -374 195 -340
<< viali >>
rect -19 238 19 272
rect -81 -188 -47 188
rect 47 -188 81 188
rect -19 -272 19 -238
<< metal1 >>
rect -31 272 31 278
rect -31 238 -19 272
rect 19 238 31 272
rect -31 232 31 238
rect -87 188 -41 200
rect -87 -188 -81 188
rect -47 -188 -41 188
rect -87 -200 -41 -188
rect 41 188 87 200
rect 41 -188 47 188
rect 81 -188 87 188
rect 41 -200 87 -188
rect -31 -238 31 -232
rect -31 -272 -19 -238
rect 19 -272 31 -238
rect -31 -278 31 -272
<< properties >>
string FIXED_BBOX -178 -357 178 357
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
