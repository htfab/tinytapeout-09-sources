magic
tech sky130A
magscale 1 2
timestamp 1730191042
<< error_p >>
rect -29 345 29 351
rect -29 311 -17 345
rect -29 305 29 311
<< nwell >>
rect -109 -398 109 364
<< pmos >>
rect -15 -336 15 264
<< pdiff >>
rect -73 252 -15 264
rect -73 -324 -61 252
rect -27 -324 -15 252
rect -73 -336 -15 -324
rect 15 252 73 264
rect 15 -324 27 252
rect 61 -324 73 252
rect 15 -336 73 -324
<< pdiffc >>
rect -61 -324 -27 252
rect 27 -324 61 252
<< poly >>
rect -33 345 33 361
rect -33 311 -17 345
rect 17 311 33 345
rect -33 295 33 311
rect -15 264 15 295
rect -15 -362 15 -336
<< polycont >>
rect -17 311 17 345
<< locali >>
rect -33 311 -17 345
rect 17 311 33 345
rect -61 252 -27 268
rect -61 -340 -27 -324
rect 27 252 61 268
rect 27 -340 61 -324
<< viali >>
rect -17 311 17 345
rect -61 -324 -27 252
rect 27 -324 61 252
<< metal1 >>
rect -29 345 29 351
rect -29 311 -17 345
rect 17 311 29 345
rect -29 305 29 311
rect -67 252 -21 264
rect -67 -324 -61 252
rect -27 -324 -21 252
rect -67 -336 -21 -324
rect 21 252 67 264
rect 21 -324 27 252
rect 61 -324 67 252
rect 21 -336 67 -324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
