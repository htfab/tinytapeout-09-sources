magic
tech sky130A
magscale 1 2
timestamp 1730925979
<< error_p >>
rect 19 381 77 387
rect 19 347 31 381
rect 19 341 77 347
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -77 -387 -19 -381
<< nwell >>
rect -263 -519 263 519
<< pmos >>
rect -63 -300 -33 300
rect 33 -300 63 300
<< pdiff >>
rect -125 288 -63 300
rect -125 -288 -113 288
rect -79 -288 -63 288
rect -125 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 125 300
rect 63 -288 79 288
rect 113 -288 125 288
rect 63 -300 125 -288
<< pdiffc >>
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
<< nsubdiff >>
rect -227 449 -131 483
rect 131 449 227 483
rect -227 387 -193 449
rect 193 387 227 449
rect -227 -449 -193 -387
rect 193 -449 227 -387
rect -227 -483 -131 -449
rect 131 -483 227 -449
<< nsubdiffcont >>
rect -131 449 131 483
rect -227 -387 -193 387
rect 193 -387 227 387
rect -131 -483 131 -449
<< poly >>
rect 15 381 81 397
rect 15 347 31 381
rect 65 347 81 381
rect 15 331 81 347
rect -63 300 -33 326
rect 33 300 63 331
rect -63 -331 -33 -300
rect 33 -326 63 -300
rect -81 -347 -15 -331
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -81 -397 -15 -381
<< polycont >>
rect 31 347 65 381
rect -65 -381 -31 -347
<< locali >>
rect -227 449 -131 483
rect 131 449 227 483
rect -227 387 -193 449
rect 193 387 227 449
rect 15 347 31 381
rect 65 347 81 381
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect -81 -381 -65 -347
rect -31 -381 -15 -347
rect -227 -449 -193 -387
rect 193 -449 227 -387
rect -227 -483 -131 -449
rect 131 -483 227 -449
<< viali >>
rect 31 347 65 381
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect -65 -381 -31 -347
<< metal1 >>
rect 19 381 77 387
rect 19 347 31 381
rect 65 347 77 381
rect 19 341 77 347
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect -77 -347 -19 -341
rect -77 -381 -65 -347
rect -31 -381 -19 -347
rect -77 -387 -19 -381
<< properties >>
string FIXED_BBOX -210 -466 210 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
