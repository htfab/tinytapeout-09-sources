* NGSPICE file created from saff_parax.ext - technology: sky130A

.subckt saff_parax d nd clk q nq VDD VSS
X0 a_3948_n831# q.t4 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X1 nq.t1 a_4216_n928# a_3948_n831# VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X2 VSS.t7 a_2276_n1548.t4 a_2236_n1460# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 a_2560_620.t1 a_2604_1734# a_2432_2796.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X4 VDD.t15 clk.t0 a_2276_n1548.t3 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X5 a_3948_n1460# q.t5 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6 a_2276_n1548.t2 a_2432_2796.t4 a_3076_620.t0 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X7 a_4216_n928# a_2432_2796.t5 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X8 a_2748_2868# a_2276_n1548.t5 a_2432_2796.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X9 VSS.t11 clk.t1 a_2652_620.t2 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X10 VSS.t9 clk.t2 a_2652_620.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X11 a_2956_n831# a_2236_n1460# q.t1 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X12 a_2652_620.t5 d.t0 a_2560_620.t4 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X13 a_2652_620.t0 clk.t3 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X14 VDD.t5 nq.t4 a_2956_n831# VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X15 a_2560_620.t3 d.t1 a_2652_620.t4 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X16 a_2652_620.t3 d.t2 a_2560_620.t2 VSS.t24 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X17 a_3076_620.t1 a_3120_1734# a_2276_n1548.t1 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X18 a_3076_620.t4 nd.t0 a_2652_620.t8 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X19 a_2652_620.t7 nd.t1 a_3076_620.t3 VSS.t25 sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X20 a_2652_620.t6 nd.t2 a_3076_620.t2 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X21 VDD.t3 a_2276_n1548.t6 a_2236_n1460# VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X22 a_2432_2796.t3 clk.t4 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X23 nq.t2 a_2276_n1548.t7 a_3948_n1460# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X24 a_2956_n1460# a_2432_2796.t6 q.t3 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X25 a_4216_n928# a_2432_2796.t7 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X26 a_2432_2796.t1 a_2276_n1548.t8 a_2560_620.t0 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X27 a_2276_n1548.t0 a_2432_2796.t8 a_2748_2868# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X28 VDD.t19 a_2276_n1548.t9 nq.t3 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X29 q.t0 a_2236_n1460# VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X30 VSS.t22 nq.t5 a_2956_n1460# VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 q.t2 a_2432_2796.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X32 VSS.t15 a_4216_n928# nq.t0 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
R0 q.t5 q.t4 1099.21
R1 q.n3 q.t5 387.947
R2 q.n0 q.t1 84.2168
R3 q.n2 q.t3 83.9618
R4 q.n0 q.t2 83.8097
R5 q.n1 q.t0 83.7172
R6 q.n3 q.n2 4.86301
R7 q.n1 q.n0 1.72958
R8 q q.n3 0.848714
R9 q.n2 q.n1 0.00159649
R10 VDD.n60 VDD.n59 2142.35
R11 VDD.n77 VDD.n73 2142.35
R12 VDD.n29 VDD.n25 2142.35
R13 VDD.n45 VDD.n7 2142.35
R14 VDD.n137 VDD.n99 2018.82
R15 VDD.n136 VDD.n99 2018.82
R16 VDD.n128 VDD.n126 2018.82
R17 VDD.n115 VDD.n105 2018.82
R18 VDD.n120 VDD.n101 2018.82
R19 VDD.n120 VDD.n102 2018.82
R20 VDD.n63 VDD.n52 1584.71
R21 VDD.n63 VDD.n57 1584.71
R22 VDD.n88 VDD.n51 1584.71
R23 VDD.n56 VDD.n51 1584.71
R24 VDD.n70 VDD.n68 1584.71
R25 VDD.n70 VDD.n66 1584.71
R26 VDD.n16 VDD.n15 1584.71
R27 VDD.n16 VDD.n13 1584.71
R28 VDD.n22 VDD.n19 1584.71
R29 VDD.n22 VDD.n21 1584.71
R30 VDD.n10 VDD.n6 1584.71
R31 VDD.n10 VDD.n9 1584.71
R32 VDD.n132 VDD.n100 1461.18
R33 VDD.n132 VDD.n124 1461.18
R34 VDD.n109 VDD.n108 1461.18
R35 VDD.n108 VDD.n106 1461.18
R36 VDD.n137 VDD.n100 557.648
R37 VDD.n128 VDD.n100 557.648
R38 VDD.n136 VDD.n124 557.648
R39 VDD.n130 VDD.n124 557.648
R40 VDD.n113 VDD.n109 557.648
R41 VDD.n109 VDD.n101 557.648
R42 VDD.n115 VDD.n106 557.648
R43 VDD.n106 VDD.n102 557.648
R44 VDD.n89 VDD.n88 557.648
R45 VDD.n88 VDD.n87 557.648
R46 VDD.n87 VDD.n52 557.648
R47 VDD.n81 VDD.n52 557.648
R48 VDD.n81 VDD.n68 557.648
R49 VDD.n77 VDD.n68 557.648
R50 VDD.n60 VDD.n56 557.648
R51 VDD.n86 VDD.n56 557.648
R52 VDD.n86 VDD.n57 557.648
R53 VDD.n82 VDD.n57 557.648
R54 VDD.n82 VDD.n66 557.648
R55 VDD.n75 VDD.n66 557.648
R56 VDD.n27 VDD.n19 557.648
R57 VDD.n34 VDD.n19 557.648
R58 VDD.n34 VDD.n15 557.648
R59 VDD.n38 VDD.n15 557.648
R60 VDD.n38 VDD.n6 557.648
R61 VDD.n45 VDD.n6 557.648
R62 VDD.n29 VDD.n21 557.648
R63 VDD.n33 VDD.n21 557.648
R64 VDD.n33 VDD.n13 557.648
R65 VDD.n39 VDD.n13 557.648
R66 VDD.n39 VDD.n9 557.648
R67 VDD.n43 VDD.n9 557.648
R68 VDD.n74 VDD.n72 228.518
R69 VDD.n61 VDD.n48 228.518
R70 VDD.n42 VDD.n4 228.518
R71 VDD.n30 VDD.n24 228.518
R72 VDD.n135 VDD.n97 215.341
R73 VDD.n131 VDD.n125 215.341
R74 VDD.n119 VDD.n118 215.341
R75 VDD.n116 VDD.n104 215.341
R76 VDD.n127 VDD.n125 211.06
R77 VDD.n122 VDD.n121 196.281
R78 VDD.n78 VDD.n72 176.998
R79 VDD.n26 VDD.n24 176.998
R80 VDD.n79 VDD.n71 169.036
R81 VDD.n71 VDD.n65 169.036
R82 VDD.n69 VDD.n64 169.036
R83 VDD.n84 VDD.n64 169.036
R84 VDD.n58 VDD.n49 169.036
R85 VDD.n62 VDD.n58 169.036
R86 VDD.n91 VDD.n48 169.036
R87 VDD.n11 VDD.n5 169.036
R88 VDD.n41 VDD.n11 169.036
R89 VDD.n36 VDD.n17 169.036
R90 VDD.n17 VDD.n12 169.036
R91 VDD.n23 VDD.n18 169.036
R92 VDD.n31 VDD.n23 169.036
R93 VDD.n47 VDD.n4 169.036
R94 VDD.n112 VDD.n104 163.294
R95 VDD.n139 VDD.n97 155.859
R96 VDD.n133 VDD.n98 155.859
R97 VDD.n134 VDD.n133 155.859
R98 VDD.n111 VDD.n103 155.859
R99 VDD.n117 VDD.n103 155.859
R100 VDD.n119 VDD.n96 155.859
R101 VDD.t14 VDD.n107 155.062
R102 VDD.n107 VDD.t0 155.062
R103 VDD.n121 VDD.t0 155.062
R104 VDD.t1 VDD.n122 155.062
R105 VDD.t1 VDD.n123 155.062
R106 VDD.t12 VDD.n123 155.062
R107 VDD.n114 VDD.n105 153.352
R108 VDD.n129 VDD.n126 153.352
R109 VDD.t4 VDD.n54 144.606
R110 VDD.t6 VDD.n54 144.606
R111 VDD.t6 VDD.n55 144.606
R112 VDD.t10 VDD.n55 144.606
R113 VDD.t10 VDD.n67 144.606
R114 VDD.t2 VDD.n67 144.606
R115 VDD.t7 VDD.n20 144.606
R116 VDD.t18 VDD.n20 144.606
R117 VDD.t18 VDD.n14 144.606
R118 VDD.t9 VDD.n14 144.606
R119 VDD.t9 VDD.n8 144.606
R120 VDD.t16 VDD.n8 144.606
R121 VDD.n59 VDD.n50 144.319
R122 VDD.n76 VDD.n73 144.319
R123 VDD.n28 VDD.n25 144.319
R124 VDD.n44 VDD.n7 144.319
R125 VDD.n131 VDD.n130 92.5005
R126 VDD.n136 VDD.n135 92.5005
R127 VDD.t1 VDD.n136 92.5005
R128 VDD.n138 VDD.n137 92.5005
R129 VDD.n137 VDD.t1 92.5005
R130 VDD.n128 VDD.n127 92.5005
R131 VDD.t12 VDD.n128 92.5005
R132 VDD.n118 VDD.n102 92.5005
R133 VDD.n102 VDD.t0 92.5005
R134 VDD.n116 VDD.n115 92.5005
R135 VDD.n115 VDD.t14 92.5005
R136 VDD.n113 VDD.n112 92.5005
R137 VDD.n110 VDD.n101 92.5005
R138 VDD.n101 VDD.t0 92.5005
R139 VDD.n75 VDD.n74 92.5005
R140 VDD.n83 VDD.n82 92.5005
R141 VDD.n82 VDD.t10 92.5005
R142 VDD.n86 VDD.n85 92.5005
R143 VDD.t6 VDD.n86 92.5005
R144 VDD.n61 VDD.n60 92.5005
R145 VDD.n60 VDD.t4 92.5005
R146 VDD.n90 VDD.n89 92.5005
R147 VDD.n87 VDD.n53 92.5005
R148 VDD.n87 VDD.t6 92.5005
R149 VDD.n81 VDD.n80 92.5005
R150 VDD.t10 VDD.n81 92.5005
R151 VDD.n78 VDD.n77 92.5005
R152 VDD.n77 VDD.t2 92.5005
R153 VDD.n43 VDD.n42 92.5005
R154 VDD.n40 VDD.n39 92.5005
R155 VDD.n39 VDD.t9 92.5005
R156 VDD.n33 VDD.n32 92.5005
R157 VDD.t18 VDD.n33 92.5005
R158 VDD.n30 VDD.n29 92.5005
R159 VDD.n29 VDD.t7 92.5005
R160 VDD.n27 VDD.n26 92.5005
R161 VDD.n35 VDD.n34 92.5005
R162 VDD.n34 VDD.t18 92.5005
R163 VDD.n38 VDD.n37 92.5005
R164 VDD.t9 VDD.n38 92.5005
R165 VDD.n46 VDD.n45 92.5005
R166 VDD.n45 VDD.t16 92.5005
R167 VDD.n95 VDD.t15 84.7512
R168 VDD.n142 VDD.t13 84.7133
R169 VDD.n1 VDD.t17 84.3878
R170 VDD.n1 VDD.t5 84.38
R171 VDD.n0 VDD.t19 84.0993
R172 VDD.n2 VDD.t11 84.0793
R173 VDD.n2 VDD.t3 83.8172
R174 VDD.n0 VDD.t8 83.8097
R175 VDD.n89 VDD.n50 82.6992
R176 VDD.n76 VDD.n75 82.6992
R177 VDD.n28 VDD.n27 82.6992
R178 VDD.n44 VDD.n43 82.6992
R179 VDD.n130 VDD.n129 81.7299
R180 VDD.n114 VDD.n113 81.7299
R181 VDD.n135 VDD.n134 59.4829
R182 VDD.n134 VDD.n131 59.4829
R183 VDD.n117 VDD.n116 59.4829
R184 VDD.n118 VDD.n117 59.4829
R185 VDD.n62 VDD.n61 59.4829
R186 VDD.n85 VDD.n62 59.4829
R187 VDD.n85 VDD.n84 59.4829
R188 VDD.n84 VDD.n83 59.4829
R189 VDD.n83 VDD.n65 59.4829
R190 VDD.n74 VDD.n65 59.4829
R191 VDD.n31 VDD.n30 59.4829
R192 VDD.n32 VDD.n31 59.4829
R193 VDD.n32 VDD.n12 59.4829
R194 VDD.n40 VDD.n12 59.4829
R195 VDD.n41 VDD.n40 59.4829
R196 VDD.n42 VDD.n41 59.4829
R197 VDD.n133 VDD.n132 18.5005
R198 VDD.n132 VDD.n123 18.5005
R199 VDD.n126 VDD.n125 18.5005
R200 VDD.n99 VDD.n97 18.5005
R201 VDD.n122 VDD.n99 18.5005
R202 VDD.n108 VDD.n103 18.5005
R203 VDD.n108 VDD.n107 18.5005
R204 VDD.n120 VDD.n119 18.5005
R205 VDD.n121 VDD.n120 18.5005
R206 VDD.n105 VDD.n104 18.5005
R207 VDD.n64 VDD.n63 16.8187
R208 VDD.n63 VDD.n55 16.8187
R209 VDD.n58 VDD.n51 16.8187
R210 VDD.n54 VDD.n51 16.8187
R211 VDD.n71 VDD.n70 16.8187
R212 VDD.n70 VDD.n67 16.8187
R213 VDD.n73 VDD.n72 16.8187
R214 VDD.n59 VDD.n48 16.8187
R215 VDD.n17 VDD.n16 16.8187
R216 VDD.n16 VDD.n14 16.8187
R217 VDD.n23 VDD.n22 16.8187
R218 VDD.n22 VDD.n20 16.8187
R219 VDD.n11 VDD.n10 16.8187
R220 VDD.n10 VDD.n8 16.8187
R221 VDD.n7 VDD.n4 16.8187
R222 VDD.n25 VDD.n24 16.8187
R223 VDD.n92 VDD.n91 10.5154
R224 VDD.n140 VDD.n139 10.4341
R225 VDD.n92 VDD.n47 10.1663
R226 VDD.n91 VDD.n90 7.9627
R227 VDD.n90 VDD.n49 7.9627
R228 VDD.n53 VDD.n49 7.9627
R229 VDD.n69 VDD.n53 7.9627
R230 VDD.n80 VDD.n69 7.9627
R231 VDD.n80 VDD.n79 7.9627
R232 VDD.n79 VDD.n78 7.9627
R233 VDD.n26 VDD.n18 7.9627
R234 VDD.n35 VDD.n18 7.9627
R235 VDD.n36 VDD.n35 7.9627
R236 VDD.n37 VDD.n36 7.9627
R237 VDD.n37 VDD.n5 7.9627
R238 VDD.n46 VDD.n5 7.9627
R239 VDD.n47 VDD.n46 7.9627
R240 VDD.n95 VDD.n94 7.51118
R241 VDD.n139 VDD.n138 7.43579
R242 VDD.n138 VDD.n98 7.43579
R243 VDD.n127 VDD.n98 7.43579
R244 VDD.n112 VDD.n111 7.43579
R245 VDD.n111 VDD.n110 7.43579
R246 VDD.n110 VDD.n96 7.43579
R247 VDD.n129 VDD.t12 7.02738
R248 VDD.t14 VDD.n114 7.02738
R249 VDD.t2 VDD.n76 6.23219
R250 VDD.t4 VDD.n50 6.23219
R251 VDD.t16 VDD.n44 6.23219
R252 VDD.t7 VDD.n28 6.23219
R253 VDD.n3 VDD.n2 1.67005
R254 VDD.n3 VDD.n1 1.12087
R255 VDD.n94 VDD.n0 0.877815
R256 VDD.n94 VDD.n93 0.799559
R257 VDD.n142 VDD.n141 0.478842
R258 VDD.n141 VDD.n95 0.357554
R259 VDD.n141 VDD.n140 0.258833
R260 VDD.n93 VDD.n92 0.11675
R261 VDD.n140 VDD.n96 0.0946176
R262 VDD VDD.n142 0.0685693
R263 VDD.n93 VDD.n3 0.00386021
R264 nq.t4 nq.t5 1099.21
R265 nq.n0 nq.t4 728.907
R266 nq.n0 nq.t1 84.2168
R267 nq.n1 nq.t2 83.9797
R268 nq.n0 nq.t3 83.8097
R269 nq.n2 nq.t0 83.7196
R270 nq nq.n2 5.63264
R271 nq.n1 nq.n0 1.54704
R272 nq.n2 nq.n1 0.00170192
R273 a_2276_n1548.t9 a_2276_n1548.t7 1108.76
R274 a_2276_n1548.t6 a_2276_n1548.t4 1099.21
R275 a_2276_n1548.n3 a_2276_n1548.t6 736.819
R276 a_2276_n1548.n0 a_2276_n1548.t9 733.443
R277 a_2276_n1548.n2 a_2276_n1548.t5 717.534
R278 a_2276_n1548.n2 a_2276_n1548.t8 703.038
R279 a_2276_n1548.n4 a_2276_n1548.t3 83.9972
R280 a_2276_n1548.t0 a_2276_n1548.n4 83.8686
R281 a_2276_n1548.n1 a_2276_n1548.t1 34.2712
R282 a_2276_n1548.n1 a_2276_n1548.t2 31.2054
R283 a_2276_n1548.n0 a_2276_n1548.n3 5.67823
R284 a_2276_n1548.n3 a_2276_n1548.n2 4.5005
R285 a_2276_n1548.n0 a_2276_n1548.n1 0.80635
R286 a_2276_n1548.n4 a_2276_n1548.n0 0.780005
R287 VSS.n84 VSS.n24 2.28491e+06
R288 VSS.n136 VSS.n24 35636.1
R289 VSS.n136 VSS.n135 32757.9
R290 VSS.n111 VSS.n61 17981.1
R291 VSS.n51 VSS.n47 5203.12
R292 VSS.n60 VSS.n47 5203.12
R293 VSS.n51 VSS.n48 5203.12
R294 VSS.n60 VSS.n48 5203.12
R295 VSS.n8 VSS.n6 4623.71
R296 VSS.n153 VSS.n6 4623.71
R297 VSS.n23 VSS.n21 4623.71
R298 VSS.n23 VSS.n22 4623.71
R299 VSS.n147 VSS.n15 3766.18
R300 VSS.n143 VSS.n15 3766.18
R301 VSS.n147 VSS.n16 3766.18
R302 VSS.n143 VSS.n16 3766.18
R303 VSS.n151 VSS.n10 3766.18
R304 VSS.n151 VSS.n11 3766.18
R305 VSS.n10 VSS.n9 3766.18
R306 VSS.n11 VSS.n9 3766.18
R307 VSS.n20 VSS.n19 3128.82
R308 VSS.n19 VSS.n7 3128.82
R309 VSS.n115 VSS.n44 2306.06
R310 VSS.n116 VSS.n44 2306.06
R311 VSS.n134 VSS.n25 2306.06
R312 VSS.n134 VSS.n26 2306.06
R313 VSS.n86 VSS.n83 2306.06
R314 VSS.n109 VSS.n62 2306.06
R315 VSS.n109 VSS.n63 2306.06
R316 VSS.n87 VSS.n83 2306.06
R317 VSS.n20 VSS.n8 1494.88
R318 VSS.n21 VSS.n20 1494.88
R319 VSS.n153 VSS.n7 1494.88
R320 VSS.n22 VSS.n7 1494.88
R321 VSS.n36 VSS.n35 1390.59
R322 VSS.n35 VSS.n31 1390.59
R323 VSS.n37 VSS.n34 1390.59
R324 VSS.n37 VSS.n30 1390.59
R325 VSS.n118 VSS.n40 1390.59
R326 VSS.n118 VSS.n42 1390.59
R327 VSS.n73 VSS.n72 1390.59
R328 VSS.n72 VSS.n68 1390.59
R329 VSS.n74 VSS.n71 1390.59
R330 VSS.n74 VSS.n67 1390.59
R331 VSS.n80 VSS.n77 1390.59
R332 VSS.n80 VSS.n79 1390.59
R333 VSS.n115 VSS.n40 915.471
R334 VSS.n123 VSS.n40 915.471
R335 VSS.n123 VSS.n34 915.471
R336 VSS.n128 VSS.n34 915.471
R337 VSS.n128 VSS.n36 915.471
R338 VSS.n36 VSS.n25 915.471
R339 VSS.n116 VSS.n42 915.471
R340 VSS.n122 VSS.n42 915.471
R341 VSS.n122 VSS.n30 915.471
R342 VSS.n129 VSS.n30 915.471
R343 VSS.n129 VSS.n31 915.471
R344 VSS.n31 VSS.n26 915.471
R345 VSS.n86 VSS.n77 915.471
R346 VSS.n92 VSS.n77 915.471
R347 VSS.n92 VSS.n71 915.471
R348 VSS.n97 VSS.n71 915.471
R349 VSS.n97 VSS.n73 915.471
R350 VSS.n73 VSS.n62 915.471
R351 VSS.n87 VSS.n79 915.471
R352 VSS.n91 VSS.n79 915.471
R353 VSS.n91 VSS.n67 915.471
R354 VSS.n98 VSS.n67 915.471
R355 VSS.n98 VSS.n68 915.471
R356 VSS.n68 VSS.n63 915.471
R357 VSS.n111 VSS.n110 733.333
R358 VSS.n112 VSS.n111 733.333
R359 VSS.n144 VSS.n136 651.73
R360 VSS.t17 VSS.n84 643.705
R361 VSS.t17 VSS.n78 643.705
R362 VSS.t14 VSS.n78 643.705
R363 VSS.t14 VSS.n69 643.705
R364 VSS.t5 VSS.n69 643.705
R365 VSS.t5 VSS.n70 643.705
R366 VSS.n70 VSS.t19 643.705
R367 VSS.n110 VSS.t19 643.705
R368 VSS.t21 VSS.n112 643.705
R369 VSS.t21 VSS.n41 643.705
R370 VSS.t23 VSS.n41 643.705
R371 VSS.t23 VSS.n32 643.705
R372 VSS.t2 VSS.n32 643.705
R373 VSS.t2 VSS.n33 643.705
R374 VSS.n33 VSS.t6 643.705
R375 VSS.n135 VSS.t6 643.705
R376 VSS.n50 VSS.n24 535.941
R377 VSS.n53 VSS.n52 338.072
R378 VSS.n132 VSS.n26 292.5
R379 VSS.n26 VSS.t6 292.5
R380 VSS.n130 VSS.n129 292.5
R381 VSS.n129 VSS.t2 292.5
R382 VSS.n122 VSS.n121 292.5
R383 VSS.t23 VSS.n122 292.5
R384 VSS.n117 VSS.n116 292.5
R385 VSS.n116 VSS.t21 292.5
R386 VSS.n115 VSS.n114 292.5
R387 VSS.t21 VSS.n115 292.5
R388 VSS.n124 VSS.n123 292.5
R389 VSS.n123 VSS.t23 292.5
R390 VSS.n128 VSS.n127 292.5
R391 VSS.t2 VSS.n128 292.5
R392 VSS.n27 VSS.n25 292.5
R393 VSS.n25 VSS.t6 292.5
R394 VSS.n86 VSS.n85 292.5
R395 VSS.t17 VSS.n86 292.5
R396 VSS.n93 VSS.n92 292.5
R397 VSS.n92 VSS.t14 292.5
R398 VSS.n97 VSS.n96 292.5
R399 VSS.t5 VSS.n97 292.5
R400 VSS.n64 VSS.n62 292.5
R401 VSS.n62 VSS.t19 292.5
R402 VSS.n101 VSS.n63 292.5
R403 VSS.n63 VSS.t19 292.5
R404 VSS.n99 VSS.n98 292.5
R405 VSS.n98 VSS.t5 292.5
R406 VSS.n91 VSS.n90 292.5
R407 VSS.t14 VSS.n91 292.5
R408 VSS.n88 VSS.n87 292.5
R409 VSS.n87 VSS.t17 292.5
R410 VSS.n50 VSS.t8 267.971
R411 VSS.n61 VSS.t10 267.971
R412 VSS.n17 VSS.t12 267.971
R413 VSS.t13 VSS.n144 267.971
R414 VSS.n52 VSS.n49 254.935
R415 VSS.n150 VSS.n12 244.707
R416 VSS.n142 VSS.n13 244.707
R417 VSS.n140 VSS.n139 217.287
R418 VSS.n18 VSS.n14 209.3
R419 VSS.n141 VSS.n140 203.294
R420 VSS.n18 VSS.n5 203.294
R421 VSS.n56 VSS.n12 165.648
R422 VSS.n142 VSS.n141 165.648
R423 VSS.t8 VSS.t0 158.798
R424 VSS.t0 VSS.t10 158.798
R425 VSS.n46 VSS.n45 158.798
R426 VSS.t16 VSS.t25 158.798
R427 VSS.n146 VSS.n17 158.798
R428 VSS.t24 VSS.t4 158.798
R429 VSS.n114 VSS.n113 149.835
R430 VSS.n133 VSS.n27 149.835
R431 VSS.n85 VSS.n82 149.835
R432 VSS.n108 VSS.n64 149.835
R433 VSS.n54 VSS.n9 146.25
R434 VSS.n152 VSS.n9 146.25
R435 VSS.n151 VSS.n150 146.25
R436 VSS.n152 VSS.n151 146.25
R437 VSS.n138 VSS.n16 146.25
R438 VSS.n145 VSS.n16 146.25
R439 VSS.n15 VSS.n13 146.25
R440 VSS.n145 VSS.n15 146.25
R441 VSS.n61 VSS.n46 145.565
R442 VSS.n57 VSS.n53 143.911
R443 VSS.n139 VSS.n22 117.001
R444 VSS.t4 VSS.n22 117.001
R445 VSS.n154 VSS.n153 117.001
R446 VSS.n153 VSS.t16 117.001
R447 VSS.n55 VSS.n8 117.001
R448 VSS.t16 VSS.n8 117.001
R449 VSS.n137 VSS.n21 117.001
R450 VSS.t4 VSS.n21 117.001
R451 VSS.n49 VSS.n48 117.001
R452 VSS.t0 VSS.n48 117.001
R453 VSS.n53 VSS.n47 117.001
R454 VSS.t0 VSS.n47 117.001
R455 VSS.n75 VSS.n74 117.001
R456 VSS.n74 VSS.n69 117.001
R457 VSS.n72 VSS.n65 117.001
R458 VSS.n72 VSS.n70 117.001
R459 VSS.n119 VSS.n118 117.001
R460 VSS.n118 VSS.n41 117.001
R461 VSS.n38 VSS.n37 117.001
R462 VSS.n37 VSS.n32 117.001
R463 VSS.n35 VSS.n28 117.001
R464 VSS.n35 VSS.n33 117.001
R465 VSS.n134 VSS.n133 117.001
R466 VSS.n135 VSS.n134 117.001
R467 VSS.n113 VSS.n44 117.001
R468 VSS.n112 VSS.n44 117.001
R469 VSS.n81 VSS.n80 117.001
R470 VSS.n80 VSS.n78 117.001
R471 VSS.n83 VSS.n82 117.001
R472 VSS.n84 VSS.n83 117.001
R473 VSS.n109 VSS.n108 117.001
R474 VSS.n110 VSS.n109 117.001
R475 VSS.n45 VSS.t25 109.174
R476 VSS.n146 VSS.t24 109.174
R477 VSS.n133 VSS.n132 99.7164
R478 VSS.n88 VSS.n82 99.7164
R479 VSS.n126 VSS.n28 90.3534
R480 VSS.n131 VSS.n28 90.3534
R481 VSS.n125 VSS.n38 90.3534
R482 VSS.n38 VSS.n29 90.3534
R483 VSS.n113 VSS.n43 90.3534
R484 VSS.n119 VSS.n39 90.3534
R485 VSS.n120 VSS.n119 90.3534
R486 VSS.n95 VSS.n65 90.3534
R487 VSS.n100 VSS.n65 90.3534
R488 VSS.n94 VSS.n75 90.3534
R489 VSS.n75 VSS.n66 90.3534
R490 VSS.n81 VSS.n76 90.3534
R491 VSS.n89 VSS.n81 90.3534
R492 VSS.n108 VSS.n107 90.3534
R493 VSS.n103 VSS.t20 84.2152
R494 VSS.n103 VSS.t22 84.2035
R495 VSS.n0 VSS.t3 83.8547
R496 VSS.n102 VSS.t18 83.8511
R497 VSS.n102 VSS.t15 83.7212
R498 VSS.n0 VSS.t7 83.7186
R499 VSS.t16 VSS.n152 79.399
R500 VSS.n152 VSS.t12 79.399
R501 VSS.t4 VSS.n145 79.399
R502 VSS.n145 VSS.t13 79.399
R503 VSS.n149 VSS.n13 72.6593
R504 VSS.n150 VSS.n149 72.6593
R505 VSS.n114 VSS.n39 59.4829
R506 VSS.n124 VSS.n39 59.4829
R507 VSS.n125 VSS.n124 59.4829
R508 VSS.n127 VSS.n125 59.4829
R509 VSS.n127 VSS.n126 59.4829
R510 VSS.n126 VSS.n27 59.4829
R511 VSS.n85 VSS.n76 59.4829
R512 VSS.n93 VSS.n76 59.4829
R513 VSS.n94 VSS.n93 59.4829
R514 VSS.n96 VSS.n94 59.4829
R515 VSS.n96 VSS.n95 59.4829
R516 VSS.n95 VSS.n64 59.4829
R517 VSS.n58 VSS.n4 56.6562
R518 VSS.n148 VSS.n11 53.1823
R519 VSS.n17 VSS.n11 53.1823
R520 VSS.n12 VSS.n10 53.1823
R521 VSS.n45 VSS.n10 53.1823
R522 VSS.n143 VSS.n142 53.1823
R523 VSS.n144 VSS.n143 53.1823
R524 VSS.n148 VSS.n147 53.1823
R525 VSS.n147 VSS.n146 53.1823
R526 VSS.n59 VSS.n57 50.7808
R527 VSS.n148 VSS.n14 49.3297
R528 VSS.n149 VSS.n148 44.9974
R529 VSS.n19 VSS.n18 41.7862
R530 VSS.n19 VSS.n17 41.7862
R531 VSS.n140 VSS.n23 41.7862
R532 VSS.n144 VSS.n23 41.7862
R533 VSS.n58 VSS.n6 41.7862
R534 VSS.n46 VSS.n6 41.7862
R535 VSS.n60 VSS.n59 34.4123
R536 VSS.n61 VSS.n60 34.4123
R537 VSS.n52 VSS.n51 34.4123
R538 VSS.n51 VSS.n50 34.4123
R539 VSS.n141 VSS.n138 22.0333
R540 VSS.n54 VSS.n14 20.2497
R541 VSS.n3 VSS.n2 18.8991
R542 VSS.n3 VSS.t9 17.8391
R543 VSS.n56 VSS.n55 16.9972
R544 VSS.n49 VSS.n4 16.3802
R545 VSS.n137 VSS.n14 15.2136
R546 VSS.n155 VSS.n4 14.9158
R547 VSS.n154 VSS.n5 13.9937
R548 VSS.n139 VSS.n5 13.9937
R549 VSS.n106 VSS.n43 12.542
R550 VSS.n107 VSS.n106 12.4013
R551 VSS.n57 VSS.n56 10.8023
R552 VSS.n59 VSS.n58 10.4923
R553 VSS.n117 VSS.n43 9.36346
R554 VSS.n120 VSS.n117 9.36346
R555 VSS.n121 VSS.n120 9.36346
R556 VSS.n121 VSS.n29 9.36346
R557 VSS.n130 VSS.n29 9.36346
R558 VSS.n131 VSS.n130 9.36346
R559 VSS.n132 VSS.n131 9.36346
R560 VSS.n89 VSS.n88 9.36346
R561 VSS.n90 VSS.n89 9.36346
R562 VSS.n90 VSS.n66 9.36346
R563 VSS.n99 VSS.n66 9.36346
R564 VSS.n100 VSS.n99 9.36346
R565 VSS.n101 VSS.n100 9.36346
R566 VSS.n107 VSS.n101 9.36346
R567 VSS.n55 VSS.n54 5.03657
R568 VSS.n138 VSS.n137 5.03657
R569 VSS.n157 VSS.n1 4.7915
R570 VSS.n2 VSS.t1 3.9605
R571 VSS.n2 VSS.t11 3.9605
R572 VSS.n156 VSS.n3 2.0131
R573 VSS.n155 VSS.n154 1.46491
R574 VSS.n105 VSS.n102 1.4286
R575 VSS.n104 VSS.n1 0.967966
R576 VSS.n157 VSS.n156 0.765444
R577 VSS.n1 VSS.n0 0.460321
R578 VSS.n104 VSS.n103 0.452881
R579 VSS.n156 VSS.n155 0.202674
R580 VSS.n106 VSS.n105 0.113915
R581 VSS VSS.n157 0.053625
R582 VSS.n105 VSS.n104 0.00392466
R583 a_2432_2796.t9 a_2432_2796.t6 1108.75
R584 a_2432_2796.t5 a_2432_2796.t7 1099.21
R585 a_2432_2796.n4 a_2432_2796.t5 739.183
R586 a_2432_2796.n2 a_2432_2796.t9 731.662
R587 a_2432_2796.n3 a_2432_2796.t8 717.299
R588 a_2432_2796.n3 a_2432_2796.t4 703.274
R589 a_2432_2796.t0 a_2432_2796.n0 84.1095
R590 a_2432_2796.n0 a_2432_2796.t3 83.8305
R591 a_2432_2796.n1 a_2432_2796.t1 34.2897
R592 a_2432_2796.n1 a_2432_2796.t2 31.1862
R593 a_2432_2796.n0 a_2432_2796.n4 5.938
R594 a_2432_2796.n4 a_2432_2796.n3 4.5005
R595 a_2432_2796.n2 a_2432_2796.n1 0.773225
R596 a_2432_2796.n0 a_2432_2796.n2 0.671045
R597 a_2560_620.n1 a_2560_620.n0 29.0038
R598 a_2560_620.n1 a_2560_620.t4 23.1697
R599 a_2560_620.n2 a_2560_620.n1 21.4537
R600 a_2560_620.n0 a_2560_620.t0 6.6005
R601 a_2560_620.n0 a_2560_620.t1 6.6005
R602 a_2560_620.t2 a_2560_620.n2 4.9505
R603 a_2560_620.n2 a_2560_620.t3 4.9505
R604 clk.n0 clk.t1 908.789
R605 clk.n0 clk.t2 908.789
R606 clk.n0 clk.t3 838.681
R607 clk.n1 clk.t0 721.708
R608 clk.n2 clk.t4 721.707
R609 clk.n1 clk.n0 169.52
R610 clk.n2 clk.n1 1.6691
R611 clk clk.n2 0.827943
R612 a_3076_620.n2 a_3076_620.n0 29.0022
R613 a_3076_620.t2 a_3076_620.n2 23.1697
R614 a_3076_620.n2 a_3076_620.n1 21.4537
R615 a_3076_620.n0 a_3076_620.t0 6.6005
R616 a_3076_620.n0 a_3076_620.t1 6.6005
R617 a_3076_620.n1 a_3076_620.t3 4.9505
R618 a_3076_620.n1 a_3076_620.t4 4.9505
R619 a_2652_620.n2 a_2652_620.t3 24.8011
R620 a_2652_620.n5 a_2652_620.t7 24.8011
R621 a_2652_620.t2 a_2652_620.n6 20.2978
R622 a_2652_620.n2 a_2652_620.n1 19.9537
R623 a_2652_620.n4 a_2652_620.n3 19.8511
R624 a_2652_620.n6 a_2652_620.n0 16.4403
R625 a_2652_620.n1 a_2652_620.t4 4.9505
R626 a_2652_620.n1 a_2652_620.t5 4.9505
R627 a_2652_620.n3 a_2652_620.t8 4.9505
R628 a_2652_620.n3 a_2652_620.t6 4.9505
R629 a_2652_620.n0 a_2652_620.t1 3.9605
R630 a_2652_620.n0 a_2652_620.t0 3.9605
R631 a_2652_620.n4 a_2652_620.n2 0.173577
R632 a_2652_620.n6 a_2652_620.n5 0.169303
R633 a_2652_620.n5 a_2652_620.n4 0.103064
R634 d.n1 d.t0 748.122
R635 d.n1 d.t2 748.122
R636 d.t0 d.n0 726.721
R637 d.n0 d.t2 726.721
R638 d.n0 d.t1 688.716
R639 d.n1 d.t1 678.014
R640 d d.n1 171.333
R641 nd.n2 nd.t2 678.014
R642 nd.n0 nd.t1 678.014
R643 nd.n1 nd.t0 678.014
R644 nd.n3 nd.n2 161.514
R645 nd.n3 nd.n0 161.514
R646 nd.n1 nd.n0 70.1096
R647 nd.n2 nd.n1 70.1096
R648 nd nd.n3 9.89419
C0 q a_2956_n831# 0.481121f
C1 a_3948_n831# nq 0.510191f
C2 VDD a_3120_1734# 0.002811f
C3 a_3948_n831# VDD 0.976456f
C4 a_4216_n928# a_2236_n1460# 0.012927f
C5 clk a_2604_1734# 2.72e-19
C6 nq nd 0.080051f
C7 d clk 0.14213f
C8 nq a_3948_n1460# 0.16713f
C9 nd VDD 0.16928f
C10 VDD a_3948_n1460# 0.012779f
C11 VDD a_2748_2868# 0.652526f
C12 nq a_2956_n831# 0.040726f
C13 VDD a_2956_n831# 0.977045f
C14 clk a_3120_1734# 8.11e-19
C15 a_3948_n831# clk 7.87e-20
C16 a_3948_n831# a_4216_n928# 0.0543f
C17 a_2956_n1460# a_2236_n1460# 0.01066f
C18 d a_2604_1734# 0.010943f
C19 nq q 0.191674f
C20 q VDD 1.44288f
C21 nd clk 0.329921f
C22 nd a_4216_n928# 4.07e-19
C23 a_3948_n1460# a_4216_n928# 0.010201f
C24 clk a_2748_2868# 0.09796f
C25 a_3120_1734# a_2604_1734# 0.002276f
C26 d a_3120_1734# 3.14e-19
C27 nd d 0.019276f
C28 q clk 0.001201f
C29 nq VDD 1.95949f
C30 q a_4216_n928# 0.040158f
C31 a_2956_n831# a_2236_n1460# 0.054279f
C32 d a_2748_2868# 0.003029f
C33 nd a_3120_1734# 0.005599f
C34 a_2956_n1460# a_2956_n831# 0.016408f
C35 q a_2236_n1460# 0.304142f
C36 a_3948_n831# a_3948_n1460# 0.016741f
C37 q d 3.69e-19
C38 nq clk 1.51e-19
C39 clk VDD 1.30375f
C40 nq a_4216_n928# 0.333395f
C41 q a_2956_n1460# 0.202483f
C42 VDD a_4216_n928# 1.13387f
C43 a_3120_1734# a_2748_2868# 0.001636f
C44 nd a_2956_n831# 8.23e-19
C45 a_3948_n831# q 0.037973f
C46 nq a_2236_n1460# 0.041577f
C47 VDD a_2236_n1460# 1.13852f
C48 VDD a_2604_1734# 0.002621f
C49 q nd 8.65e-20
C50 d VDD 0.152321f
C51 q a_3948_n1460# 0.031858f
C52 nq a_2956_n1460# 0.029749f
C53 VDD a_2956_n1460# 0.012838f
C54 nq VSS 1.59236f
C55 q VSS 2.06192f
C56 nd VSS 2.26567f
C57 d VSS 1.67945f
C58 clk VSS 1.58578f
C59 VDD VSS 21.938858f
C60 a_3948_n1460# VSS 0.425459f
C61 a_2956_n1460# VSS 0.425923f
C62 a_4216_n928# VSS 1.20677f
C63 a_3948_n831# VSS 0.05923f
C64 a_2956_n831# VSS 0.059068f
C65 a_2236_n1460# VSS 1.27378f
C66 a_3120_1734# VSS 0.183158f
C67 a_2604_1734# VSS 0.177872f
C68 a_2748_2868# VSS 0.076125f
C69 a_2652_620.t1 VSS 0.069266f
C70 a_2652_620.t0 VSS 0.069266f
C71 a_2652_620.n0 VSS 0.195611f
C72 a_2652_620.t4 VSS 0.055413f
C73 a_2652_620.t5 VSS 0.055413f
C74 a_2652_620.n1 VSS 0.146838f
C75 a_2652_620.t3 VSS 0.204997f
C76 a_2652_620.n2 VSS 0.916463f
C77 a_2652_620.t8 VSS 0.055413f
C78 a_2652_620.t6 VSS 0.055413f
C79 a_2652_620.n3 VSS 0.144904f
C80 a_2652_620.n4 VSS 0.50489f
C81 a_2652_620.t7 VSS 0.204997f
C82 a_2652_620.n5 VSS 0.538261f
C83 a_2652_620.n6 VSS 1.01603f
C84 a_2652_620.t2 VSS 0.266826f
C85 a_3076_620.t0 VSS 0.047397f
C86 a_3076_620.t1 VSS 0.047397f
C87 a_3076_620.n0 VSS 0.169349f
C88 a_3076_620.t3 VSS 0.063197f
C89 a_3076_620.t4 VSS 0.063197f
C90 a_3076_620.n1 VSS 0.207256f
C91 a_3076_620.n2 VSS 1.59121f
C92 a_3076_620.t2 VSS 0.210997f
C93 a_2560_620.t3 VSS 0.055301f
C94 a_2560_620.t0 VSS 0.041476f
C95 a_2560_620.t1 VSS 0.041476f
C96 a_2560_620.n0 VSS 0.148171f
C97 a_2560_620.t4 VSS 0.184637f
C98 a_2560_620.n1 VSS 1.39227f
C99 a_2560_620.n2 VSS 0.181364f
C100 a_2560_620.t2 VSS 0.055301f
C101 a_2432_2796.n0 VSS 0.908188f
C102 a_2432_2796.t2 VSS 0.179273f
C103 a_2432_2796.t1 VSS 0.221208f
C104 a_2432_2796.n1 VSS 0.977583f
C105 a_2432_2796.t6 VSS 0.301253f
C106 a_2432_2796.t9 VSS 0.217057f
C107 a_2432_2796.n2 VSS 1.36434f
C108 a_2432_2796.t7 VSS 0.199551f
C109 a_2432_2796.t5 VSS 0.176999f
C110 a_2432_2796.t8 VSS 0.085404f
C111 a_2432_2796.t4 VSS 0.084801f
C112 a_2432_2796.n3 VSS 0.23665f
C113 a_2432_2796.n4 VSS 1.99305f
C114 a_2432_2796.t3 VSS 0.176874f
C115 a_2432_2796.t0 VSS 0.177766f
C116 a_2276_n1548.n0 VSS 1.56413f
C117 a_2276_n1548.t3 VSS 0.164981f
C118 a_2276_n1548.t2 VSS 0.167298f
C119 a_2276_n1548.t1 VSS 0.206126f
C120 a_2276_n1548.n1 VSS 0.876206f
C121 a_2276_n1548.t7 VSS 0.281767f
C122 a_2276_n1548.t9 VSS 0.204699f
C123 a_2276_n1548.t4 VSS 0.186075f
C124 a_2276_n1548.t6 VSS 0.159193f
C125 a_2276_n1548.t5 VSS 0.079666f
C126 a_2276_n1548.t8 VSS 0.079031f
C127 a_2276_n1548.n2 VSS 0.22068f
C128 a_2276_n1548.n3 VSS 1.51054f
C129 a_2276_n1548.n4 VSS 0.434594f
C130 a_2276_n1548.t0 VSS 0.165013f
C131 VDD.t13 VSS 0.023462f
C132 VDD.t15 VSS 0.023466f
C133 VDD.t19 VSS 0.023017f
C134 VDD.t8 VSS 0.023003f
C135 VDD.n0 VSS 0.039437f
C136 VDD.t17 VSS 0.02305f
C137 VDD.t5 VSS 0.023049f
C138 VDD.n1 VSS 0.036453f
C139 VDD.t11 VSS 0.023017f
C140 VDD.t3 VSS 0.023004f
C141 VDD.n2 VSS 0.099587f
C142 VDD.n3 VSS 0.156689f
C143 VDD.n4 VSS 0.012964f
C144 VDD.n5 VSS 0.034206f
C145 VDD.n6 VSS 0.009313f
C146 VDD.n7 VSS 0.102893f
C147 VDD.n8 VSS 0.117448f
C148 VDD.n9 VSS 0.009313f
C149 VDD.n10 VSS 0.010932f
C150 VDD.n11 VSS 0.010932f
C151 VDD.n12 VSS 0.009313f
C152 VDD.n13 VSS 0.009313f
C153 VDD.n14 VSS 0.117448f
C154 VDD.n15 VSS 0.009313f
C155 VDD.n16 VSS 0.010932f
C156 VDD.n17 VSS 0.010932f
C157 VDD.n18 VSS 0.034206f
C158 VDD.n19 VSS 0.009313f
C159 VDD.n20 VSS 0.117448f
C160 VDD.n21 VSS 0.009313f
C161 VDD.n22 VSS 0.010932f
C162 VDD.n23 VSS 0.010932f
C163 VDD.n24 VSS 0.013726f
C164 VDD.n25 VSS 0.102893f
C165 VDD.n26 VSS 0.044919f
C166 VDD.n27 VSS 0.009619f
C167 VDD.t7 VSS 0.127671f
C168 VDD.n29 VSS 0.009619f
C169 VDD.n30 VSS 0.009619f
C170 VDD.n31 VSS 0.009313f
C171 VDD.n32 VSS 0.003847f
C172 VDD.n33 VSS 0.003847f
C173 VDD.t18 VSS 0.117448f
C174 VDD.n34 VSS 0.003847f
C175 VDD.n35 VSS 0.02874f
C176 VDD.n36 VSS 0.034206f
C177 VDD.n37 VSS 0.02874f
C178 VDD.n38 VSS 0.003847f
C179 VDD.t9 VSS 0.117448f
C180 VDD.n39 VSS 0.003847f
C181 VDD.n40 VSS 0.003847f
C182 VDD.n41 VSS 0.009313f
C183 VDD.n42 VSS 0.009619f
C184 VDD.n43 VSS 0.009619f
C185 VDD.t16 VSS 0.127671f
C186 VDD.n45 VSS 0.009619f
C187 VDD.n46 VSS 0.02874f
C188 VDD.n47 VSS 0.03434f
C189 VDD.n48 VSS 0.012964f
C190 VDD.n49 VSS 0.034206f
C191 VDD.n51 VSS 0.010932f
C192 VDD.n52 VSS 0.009313f
C193 VDD.n53 VSS 0.02874f
C194 VDD.n54 VSS 0.117448f
C195 VDD.n55 VSS 0.117448f
C196 VDD.n56 VSS 0.009313f
C197 VDD.n57 VSS 0.009313f
C198 VDD.n58 VSS 0.010932f
C199 VDD.n59 VSS 0.102893f
C200 VDD.t4 VSS 0.127671f
C201 VDD.n60 VSS 0.009619f
C202 VDD.n61 VSS 0.009619f
C203 VDD.n62 VSS 0.009313f
C204 VDD.n63 VSS 0.010932f
C205 VDD.n64 VSS 0.010932f
C206 VDD.n65 VSS 0.009313f
C207 VDD.n66 VSS 0.009313f
C208 VDD.n67 VSS 0.117448f
C209 VDD.n68 VSS 0.009313f
C210 VDD.n69 VSS 0.034206f
C211 VDD.n70 VSS 0.010932f
C212 VDD.n71 VSS 0.010932f
C213 VDD.n72 VSS 0.01374f
C214 VDD.n73 VSS 0.102893f
C215 VDD.n74 VSS 0.009619f
C216 VDD.n75 VSS 0.009619f
C217 VDD.t2 VSS 0.127671f
C218 VDD.n77 VSS 0.009619f
C219 VDD.n78 VSS 0.04522f
C220 VDD.n79 VSS 0.034206f
C221 VDD.n80 VSS 0.02874f
C222 VDD.n81 VSS 0.003847f
C223 VDD.t10 VSS 0.117448f
C224 VDD.n82 VSS 0.003847f
C225 VDD.n83 VSS 0.003847f
C226 VDD.n84 VSS 0.009313f
C227 VDD.n85 VSS 0.003847f
C228 VDD.n86 VSS 0.003847f
C229 VDD.t6 VSS 0.117448f
C230 VDD.n87 VSS 0.003847f
C231 VDD.n88 VSS 0.009313f
C232 VDD.n89 VSS 0.009619f
C233 VDD.n90 VSS 0.02874f
C234 VDD.n91 VSS 0.034813f
C235 VDD.n92 VSS 0.028064f
C236 VDD.n93 VSS 0.07952f
C237 VDD.n94 VSS 0.27271f
C238 VDD.n95 VSS 0.247718f
C239 VDD.n96 VSS 0.020623f
C240 VDD.n97 VSS 0.012118f
C241 VDD.n98 VSS 0.035816f
C242 VDD.n99 VSS 0.014156f
C243 VDD.n100 VSS 0.008887f
C244 VDD.t0 VSS 0.109527f
C245 VDD.n101 VSS 0.009187f
C246 VDD.n102 VSS 0.009187f
C247 VDD.n103 VSS 0.01008f
C248 VDD.n104 VSS 0.01292f
C249 VDD.n105 VSS 0.095907f
C250 VDD.n106 VSS 0.008887f
C251 VDD.n107 VSS 0.109527f
C252 VDD.n108 VSS 0.01008f
C253 VDD.n109 VSS 0.008887f
C254 VDD.n110 VSS 0.030776f
C255 VDD.n111 VSS 0.035816f
C256 VDD.n112 VSS 0.047579f
C257 VDD.n113 VSS 0.009187f
C258 VDD.t14 VSS 0.119281f
C259 VDD.n115 VSS 0.009187f
C260 VDD.n116 VSS 0.009187f
C261 VDD.n117 VSS 0.008887f
C262 VDD.n118 VSS 0.009187f
C263 VDD.n119 VSS 0.012118f
C264 VDD.n120 VSS 0.014156f
C265 VDD.n121 VSS 0.124085f
C266 VDD.n122 VSS 0.124085f
C267 VDD.n123 VSS 0.109527f
C268 VDD.n124 VSS 0.008887f
C269 VDD.n125 VSS 0.014015f
C270 VDD.n126 VSS 0.095907f
C271 VDD.n127 VSS 0.025008f
C272 VDD.n128 VSS 0.009187f
C273 VDD.t12 VSS 0.119281f
C274 VDD.n130 VSS 0.009187f
C275 VDD.n131 VSS 0.009187f
C276 VDD.n132 VSS 0.01008f
C277 VDD.n133 VSS 0.01008f
C278 VDD.n134 VSS 0.008887f
C279 VDD.n135 VSS 0.009187f
C280 VDD.n136 VSS 0.009187f
C281 VDD.t1 VSS 0.109527f
C282 VDD.n137 VSS 0.009187f
C283 VDD.n138 VSS 0.030776f
C284 VDD.n139 VSS 0.03773f
C285 VDD.n140 VSS 0.017419f
C286 VDD.n141 VSS 0.097644f
C287 VDD.n142 VSS 0.120072f
.ends

