magic
tech sky130A
timestamp 1730931062
<< locali >>
rect -170 -330 -120 -320
rect -170 -380 300 -330
rect 460 -420 710 -370
rect -360 -950 -350 -860
rect -120 -1150 960 -1100
<< viali >>
rect -500 -310 -470 -280
rect -450 -310 -420 -280
rect -400 -310 -370 -280
rect -350 -310 -320 -280
rect -300 -310 -270 -280
rect -250 -310 -220 -280
rect 440 -370 470 -340
rect 490 -370 520 -340
rect 540 -370 570 -340
rect 590 -370 620 -340
rect 640 -370 670 -340
rect 690 -370 720 -340
rect 1470 -1090 1500 -1060
rect 1520 -1090 1550 -1060
rect 1570 -1090 1600 -1060
rect 1620 -1090 1650 -1060
rect 1670 -1090 1700 -1060
rect 1720 -1090 1750 -1060
rect -500 -1140 -470 -1110
rect -450 -1140 -420 -1110
rect -400 -1140 -370 -1110
rect -350 -1140 -320 -1110
rect -300 -1140 -270 -1110
rect -250 -1140 -220 -1110
<< metal1 >>
rect -600 -250 1100 -200
rect -600 -370 -550 -250
rect -510 -280 -210 -270
rect -510 -310 -500 -280
rect -470 -310 -450 -280
rect -420 -310 -400 -280
rect -370 -310 -350 -280
rect -320 -310 -300 -280
rect -270 -310 -250 -280
rect -220 -310 -210 -280
rect -510 -320 -210 -310
rect 430 -340 730 -330
rect 430 -370 440 -340
rect 470 -370 490 -340
rect 520 -370 540 -340
rect 570 -370 590 -340
rect 620 -370 640 -340
rect 670 -370 690 -340
rect 720 -370 730 -340
rect 430 -380 730 -370
rect -120 -610 300 -600
rect -120 -640 110 -610
rect 140 -640 300 -610
rect -120 -650 300 -640
rect -150 -750 -120 -700
rect 300 -750 350 -700
rect 1460 -1060 1760 -1050
rect 1460 -1090 1470 -1060
rect 1500 -1090 1520 -1060
rect 1550 -1090 1570 -1060
rect 1600 -1090 1620 -1060
rect 1650 -1090 1670 -1060
rect 1700 -1090 1720 -1060
rect 1750 -1090 1760 -1060
rect 1460 -1100 1760 -1090
rect -510 -1110 -210 -1100
rect -510 -1140 -500 -1110
rect -470 -1140 -450 -1110
rect -420 -1140 -400 -1110
rect -370 -1140 -350 -1110
rect -320 -1140 -300 -1110
rect -270 -1140 -250 -1110
rect -220 -1140 -210 -1110
rect -510 -1150 -210 -1140
<< via1 >>
rect -500 -310 -470 -280
rect -450 -310 -420 -280
rect -400 -310 -370 -280
rect -350 -310 -320 -280
rect -300 -310 -270 -280
rect -250 -310 -220 -280
rect 440 -370 470 -340
rect 490 -370 520 -340
rect 540 -370 570 -340
rect 590 -370 620 -340
rect 640 -370 670 -340
rect 690 -370 720 -340
rect 110 -640 140 -610
rect -370 -740 -340 -710
rect 850 -740 880 -710
rect 1470 -1090 1500 -1060
rect 1520 -1090 1550 -1060
rect 1570 -1090 1600 -1060
rect 1620 -1090 1650 -1060
rect 1670 -1090 1700 -1060
rect 1720 -1090 1750 -1060
rect -500 -1140 -470 -1110
rect -450 -1140 -420 -1110
rect -400 -1140 -370 -1110
rect -350 -1140 -320 -1110
rect -300 -1140 -270 -1110
rect -250 -1140 -220 -1110
<< metal2 >>
rect -510 -280 -210 -270
rect -510 -310 -500 -280
rect -470 -310 -450 -280
rect -420 -310 -400 -280
rect -370 -310 -350 -280
rect -320 -310 -300 -280
rect -270 -310 -250 -280
rect -220 -310 -210 -280
rect -510 -320 -210 -310
rect -50 -700 0 -50
rect 100 -610 150 -50
rect 430 -340 730 -330
rect 430 -370 440 -340
rect 470 -370 490 -340
rect 520 -370 540 -340
rect 570 -370 590 -340
rect 620 -370 640 -340
rect 670 -370 690 -340
rect 720 -370 730 -340
rect 430 -380 730 -370
rect 100 -640 110 -610
rect 140 -640 150 -610
rect 100 -650 150 -640
rect 2500 -650 2600 -550
rect -380 -710 890 -700
rect -380 -740 -370 -710
rect -340 -740 850 -710
rect 880 -740 890 -710
rect -380 -750 890 -740
rect 2500 -900 2600 -800
rect 1460 -1060 1760 -1050
rect 1460 -1090 1470 -1060
rect 1500 -1090 1520 -1060
rect 1550 -1090 1570 -1060
rect 1600 -1090 1620 -1060
rect 1650 -1090 1670 -1060
rect 1700 -1090 1720 -1060
rect 1750 -1090 1760 -1060
rect 1460 -1100 1760 -1090
rect -510 -1110 -210 -1100
rect -510 -1140 -500 -1110
rect -470 -1140 -450 -1110
rect -420 -1140 -400 -1110
rect -370 -1140 -350 -1110
rect -320 -1140 -300 -1110
rect -270 -1140 -250 -1110
rect -220 -1140 -210 -1110
rect -510 -1150 -210 -1140
<< via2 >>
rect -500 -310 -470 -280
rect -450 -310 -420 -280
rect -400 -310 -370 -280
rect -350 -310 -320 -280
rect -300 -310 -270 -280
rect -250 -310 -220 -280
rect 440 -370 470 -340
rect 490 -370 520 -340
rect 540 -370 570 -340
rect 590 -370 620 -340
rect 640 -370 670 -340
rect 690 -370 720 -340
rect 1470 -1090 1500 -1060
rect 1520 -1090 1550 -1060
rect 1570 -1090 1600 -1060
rect 1620 -1090 1650 -1060
rect 1670 -1090 1700 -1060
rect 1720 -1090 1750 -1060
rect -500 -1140 -470 -1110
rect -450 -1140 -420 -1110
rect -400 -1140 -370 -1110
rect -350 -1140 -320 -1110
rect -300 -1140 -270 -1110
rect -250 -1140 -220 -1110
<< metal3 >>
rect -530 -250 -210 -220
rect -530 -310 -500 -250
rect -450 -280 -400 -250
rect -350 -280 -300 -250
rect -250 -280 -210 -250
rect -470 -310 -450 -300
rect -420 -310 -400 -280
rect -370 -310 -350 -300
rect -320 -310 -300 -280
rect -270 -310 -250 -300
rect -220 -310 -210 -280
rect -530 -320 -210 -310
rect 430 -250 730 -220
rect 430 -300 450 -250
rect 500 -300 550 -250
rect 600 -300 650 -250
rect 700 -300 730 -250
rect 430 -340 730 -300
rect 430 -370 440 -340
rect 470 -370 490 -340
rect 520 -370 540 -340
rect 570 -370 590 -340
rect 620 -370 640 -340
rect 670 -370 690 -340
rect 720 -370 730 -340
rect 430 -380 730 -370
rect 1460 -1060 1760 -1050
rect 1460 -1090 1470 -1060
rect 1500 -1090 1520 -1060
rect 1550 -1090 1570 -1060
rect 1600 -1090 1620 -1060
rect 1650 -1090 1670 -1060
rect 1700 -1090 1720 -1060
rect 1750 -1090 1760 -1060
rect 1460 -1100 1760 -1090
rect -510 -1110 -210 -1100
rect -510 -1140 -500 -1110
rect -470 -1140 -450 -1110
rect -420 -1140 -400 -1110
rect -370 -1140 -350 -1110
rect -320 -1140 -300 -1110
rect -270 -1140 -250 -1110
rect -220 -1140 -210 -1110
rect -510 -1150 -210 -1140
rect -510 -1200 -500 -1150
rect -450 -1200 -400 -1150
rect -350 -1200 -300 -1150
rect -250 -1200 -210 -1150
rect 1460 -1150 1500 -1100
rect 1550 -1150 1600 -1100
rect 1650 -1150 1700 -1100
rect 1750 -1150 1760 -1100
rect 1460 -1170 1760 -1150
rect -510 -1220 -210 -1200
<< via3 >>
rect -500 -280 -450 -250
rect -400 -280 -350 -250
rect -300 -280 -250 -250
rect -500 -300 -470 -280
rect -470 -300 -450 -280
rect -400 -300 -370 -280
rect -370 -300 -350 -280
rect -300 -300 -270 -280
rect -270 -300 -250 -280
rect 450 -300 500 -250
rect 550 -300 600 -250
rect 650 -300 700 -250
rect -500 -1200 -450 -1150
rect -400 -1200 -350 -1150
rect -300 -1200 -250 -1150
rect 1500 -1150 1550 -1100
rect 1600 -1150 1650 -1100
rect 1700 -1150 1750 -1100
<< metal4 >>
rect -1000 -250 900 -200
rect -1000 -300 -500 -250
rect -450 -300 -400 -250
rect -350 -300 -300 -250
rect -250 -300 450 -250
rect 500 -300 550 -250
rect 600 -300 650 -250
rect 700 -300 900 -250
rect -1000 -400 900 -300
rect 1460 -1100 1800 -1050
rect -1000 -1150 1500 -1100
rect 1550 -1150 1600 -1100
rect 1650 -1150 1700 -1100
rect 1750 -1150 1800 -1100
rect -1000 -1200 -500 -1150
rect -450 -1200 -400 -1150
rect -350 -1200 -300 -1150
rect -250 -1200 1800 -1150
rect -1000 -1300 1800 -1200
use SWTCH_GATE  SWTCH_GATE_0 ~/dev/personal/chacha-silicon/tt09-analog-switch/swtch_gate_sky130nm/design/SWTCH_GATE_SKY130NM
timestamp 1730928274
transform 1 0 330 0 1 -1050
box -30 -50 2200 720
use SWTCH_TWOINV  SWTCH_TWOINV_0 ~/dev/personal/chacha-silicon/tt09-analog-switch/swtch_twoinv_sky130nm/design/SWTCH_TWOINV_SKY130NM
timestamp 1730926491
transform 1 0 410 0 1 -790
box -1010 -360 -527 520
<< labels >>
rlabel metal4 -1000 -1300 -800 -1100 1 VPWR
port 1 n
rlabel metal4 -1000 -400 -800 -200 1 VGND
port 2 n
rlabel metal1 1050 -250 1100 -200 1 CTRL
port 3 n
rlabel metal2 2500 -650 2600 -550 1 X
port 4 n
rlabel metal2 2500 -900 2600 -800 1 Y
port 5 n
rlabel metal2 100 -100 150 -50 1 Q_P
port 6 n
rlabel metal2 -50 -100 0 -50 1 Q_N
port 7 n
<< end >>
