magic
tech sky130A
magscale 1 2
timestamp 1728242959
<< viali >>
rect 66 6132 1098 6168
rect 78 -18 438 18
<< metal1 >>
rect -390 6368 1230 6400
rect -390 6236 66 6368
rect 1098 6236 1230 6368
rect -390 6168 1230 6236
rect -390 6132 66 6168
rect 1098 6132 1230 6168
rect -390 6110 1230 6132
rect -182 6022 1048 6082
rect -182 1946 -118 6022
rect 170 5978 226 5984
rect 170 4402 226 4408
rect 362 5978 418 5984
rect 362 4402 418 4408
rect 554 5978 610 5984
rect 554 4402 610 4408
rect 746 5978 802 5984
rect 746 4402 802 4408
rect 938 5978 994 5984
rect 938 4402 994 4408
rect 74 3364 130 3370
rect 74 1984 130 1990
rect 266 3364 322 3370
rect 266 1984 322 1990
rect 458 3364 514 3370
rect 458 1984 514 1990
rect 650 3364 706 3370
rect 650 1984 706 1990
rect 842 3364 898 3370
rect 842 1984 898 1990
rect 1034 3364 1090 3370
rect 1034 1984 1090 1990
rect -182 1886 960 1946
rect -182 1810 298 1886
rect -390 1530 298 1810
rect -182 1386 298 1530
rect 710 1730 1210 1750
rect 710 1590 730 1730
rect 1190 1590 1210 1730
rect -182 128 -118 1386
rect 180 1350 240 1358
rect 180 942 184 1350
rect 236 942 240 1350
rect 180 934 240 942
rect 372 1350 432 1358
rect 372 942 376 1350
rect 428 942 432 1350
rect 710 1220 1210 1590
rect 372 934 432 942
rect 84 572 144 580
rect 84 164 88 572
rect 140 164 144 572
rect 84 156 144 164
rect 276 572 336 580
rect 276 164 280 572
rect 332 164 336 572
rect 276 156 336 164
rect -182 68 394 128
rect -390 18 580 40
rect -390 -18 78 18
rect 438 -18 580 18
rect -390 -82 580 -18
rect -390 -210 0 -82
rect 520 -210 580 -82
rect -390 -240 580 -210
<< via1 >>
rect 66 6236 1098 6368
rect 170 4408 226 5978
rect 362 4408 418 5978
rect 554 4408 610 5978
rect 746 4408 802 5978
rect 938 4408 994 5978
rect 74 1990 130 3364
rect 266 1990 322 3364
rect 458 1990 514 3364
rect 650 1990 706 3364
rect 842 1990 898 3364
rect 1034 1990 1090 3364
rect 730 1590 1190 1730
rect 184 942 236 1350
rect 376 942 428 1350
rect 88 164 140 572
rect 280 164 332 572
rect 0 -210 520 -82
<< metal2 >>
rect -52 6368 1218 6400
rect -52 6236 66 6368
rect 1098 6236 1218 6368
rect -52 5978 1218 6236
rect -52 4408 170 5978
rect 226 4408 362 5978
rect 418 4408 554 5978
rect 610 4408 746 5978
rect 802 4408 938 5978
rect 994 4408 1218 5978
rect -52 4402 1218 4408
rect -54 3364 1216 3370
rect -54 1990 74 3364
rect 130 1990 266 3364
rect 322 1990 458 3364
rect 514 1990 650 3364
rect 706 1990 842 3364
rect 898 1990 1034 3364
rect 1090 1990 1216 3364
rect -54 1730 1216 1990
rect -54 1590 730 1730
rect 1190 1590 1216 1730
rect -54 1568 1216 1590
rect -54 1350 570 1568
rect -54 942 184 1350
rect 236 942 376 1350
rect 428 942 570 1350
rect -54 934 570 942
rect -54 572 570 580
rect -54 164 88 572
rect 140 164 280 572
rect 332 164 570 572
rect -54 -82 570 164
rect -54 -210 0 -82
rect 520 -210 570 -82
rect -54 -238 570 -210
use sky130_fd_pr__nfet_01v8_CG2JGS  sky130_fd_pr__nfet_01v8_CG2JGS_0
timestamp 1728214159
transform 1 0 258 0 1 757
box -311 -810 311 810
use sky130_fd_pr__pfet_01v8_8DVQZL  sky130_fd_pr__pfet_01v8_8DVQZL_0
timestamp 1728214159
transform 1 0 582 0 1 3984
box -647 -2219 647 2219
<< labels >>
rlabel metal1 -390 -240 -140 10 1 VSS
rlabel metal1 -390 6110 -140 6360 1 VDD
rlabel metal1 -390 1530 -140 1780 1 in
rlabel metal1 960 1220 1210 1470 1 out
<< end >>
