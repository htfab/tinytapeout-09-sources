magic
tech sky130A
magscale 1 2
timestamp 1730889744
<< viali >>
rect 13093 27081 13127 27115
rect 13277 26945 13311 26979
rect 11253 24769 11287 24803
rect 11713 24769 11747 24803
rect 12072 24769 12106 24803
rect 14381 24769 14415 24803
rect 21373 24769 21407 24803
rect 11805 24701 11839 24735
rect 13829 24701 13863 24735
rect 11621 24633 11655 24667
rect 13185 24633 13219 24667
rect 11069 24565 11103 24599
rect 13277 24565 13311 24599
rect 14289 24565 14323 24599
rect 21189 24565 21223 24599
rect 18429 24361 18463 24395
rect 12173 24225 12207 24259
rect 18429 24225 18463 24259
rect 18521 24225 18555 24259
rect 18981 24225 19015 24259
rect 11345 24157 11379 24191
rect 11621 24157 11655 24191
rect 11805 24157 11839 24191
rect 12081 24157 12115 24191
rect 12541 24157 12575 24191
rect 14105 24157 14139 24191
rect 16313 24157 16347 24191
rect 16497 24157 16531 24191
rect 17897 24157 17931 24191
rect 18153 24157 18187 24191
rect 18613 24157 18647 24191
rect 18705 24157 18739 24191
rect 18797 24157 18831 24191
rect 21557 24157 21591 24191
rect 23029 24157 23063 24191
rect 12786 24089 12820 24123
rect 14289 24089 14323 24123
rect 18245 24089 18279 24123
rect 21290 24089 21324 24123
rect 22762 24089 22796 24123
rect 10701 24021 10735 24055
rect 11713 24021 11747 24055
rect 12449 24021 12483 24055
rect 13921 24021 13955 24055
rect 14473 24021 14507 24055
rect 16405 24021 16439 24055
rect 16773 24021 16807 24055
rect 18981 24021 19015 24055
rect 20177 24021 20211 24055
rect 21649 24021 21683 24055
rect 9413 23817 9447 23851
rect 12909 23817 12943 23851
rect 21373 23817 21407 23851
rect 8769 23749 8803 23783
rect 13645 23749 13679 23783
rect 10526 23681 10560 23715
rect 10793 23681 10827 23715
rect 10885 23681 10919 23715
rect 10977 23681 11011 23715
rect 11529 23681 11563 23715
rect 11796 23681 11830 23715
rect 13277 23681 13311 23715
rect 14565 23681 14599 23715
rect 14749 23681 14783 23715
rect 17805 23681 17839 23715
rect 18061 23681 18095 23715
rect 19073 23681 19107 23715
rect 19329 23681 19363 23715
rect 20913 23681 20947 23715
rect 21005 23681 21039 23715
rect 4905 23613 4939 23647
rect 5181 23613 5215 23647
rect 5273 23613 5307 23647
rect 5390 23613 5424 23647
rect 11161 23613 11195 23647
rect 11253 23613 11287 23647
rect 13185 23613 13219 23647
rect 13553 23613 13587 23647
rect 14289 23613 14323 23647
rect 16221 23613 16255 23647
rect 18153 23613 18187 23647
rect 20821 23613 20855 23647
rect 5549 23477 5583 23511
rect 8677 23477 8711 23511
rect 11345 23477 11379 23511
rect 13001 23477 13035 23511
rect 13737 23477 13771 23511
rect 14749 23477 14783 23511
rect 15669 23477 15703 23511
rect 16681 23477 16715 23511
rect 18797 23477 18831 23511
rect 20453 23477 20487 23511
rect 10517 23273 10551 23307
rect 11345 23273 11379 23307
rect 12173 23273 12207 23307
rect 13277 23273 13311 23307
rect 13829 23273 13863 23307
rect 18705 23273 18739 23307
rect 19257 23273 19291 23307
rect 21097 23273 21131 23307
rect 3617 23205 3651 23239
rect 12265 23205 12299 23239
rect 12541 23205 12575 23239
rect 19993 23205 20027 23239
rect 25697 23205 25731 23239
rect 4261 23137 4295 23171
rect 4629 23137 4663 23171
rect 4746 23137 4780 23171
rect 10701 23137 10735 23171
rect 11529 23137 11563 23171
rect 16497 23137 16531 23171
rect 18521 23137 18555 23171
rect 18797 23137 18831 23171
rect 21741 23137 21775 23171
rect 2237 23069 2271 23103
rect 4997 23069 5031 23103
rect 5264 23069 5298 23103
rect 7205 23069 7239 23103
rect 8953 23069 8987 23103
rect 10793 23069 10827 23103
rect 11253 23069 11287 23103
rect 11445 23063 11479 23097
rect 12449 23069 12483 23103
rect 12633 23069 12667 23103
rect 12725 23069 12759 23103
rect 12909 23069 12943 23103
rect 13277 23069 13311 23103
rect 13369 23069 13403 23103
rect 13737 23069 13771 23103
rect 13921 23069 13955 23103
rect 15413 23069 15447 23103
rect 15669 23069 15703 23103
rect 15761 23069 15795 23103
rect 16753 23069 16787 23103
rect 18705 23069 18739 23103
rect 19441 23069 19475 23103
rect 19533 23069 19567 23103
rect 19717 23069 19751 23103
rect 19809 23069 19843 23103
rect 19993 23069 20027 23103
rect 20177 23069 20211 23103
rect 20453 23069 20487 23103
rect 20913 23069 20947 23103
rect 21557 23069 21591 23103
rect 21649 23069 21683 23103
rect 21833 23069 21867 23103
rect 21925 23069 21959 23103
rect 22109 23069 22143 23103
rect 25237 23069 25271 23103
rect 25881 23069 25915 23103
rect 2504 23001 2538 23035
rect 7450 23001 7484 23035
rect 9198 23001 9232 23035
rect 11069 23001 11103 23035
rect 11161 23001 11195 23035
rect 20591 23001 20625 23035
rect 20729 23001 20763 23035
rect 20821 23001 20855 23035
rect 21373 23001 21407 23035
rect 4537 22933 4571 22967
rect 4905 22933 4939 22967
rect 6377 22933 6411 22967
rect 8585 22933 8619 22967
rect 10333 22933 10367 22967
rect 13645 22933 13679 22967
rect 14289 22933 14323 22967
rect 16405 22933 16439 22967
rect 17877 22933 17911 22967
rect 17969 22933 18003 22967
rect 19073 22933 19107 22967
rect 21189 22933 21223 22967
rect 21925 22933 21959 22967
rect 25421 22933 25455 22967
rect 2513 22729 2547 22763
rect 2881 22729 2915 22763
rect 7021 22729 7055 22763
rect 14933 22729 14967 22763
rect 15761 22729 15795 22763
rect 17877 22729 17911 22763
rect 18153 22729 18187 22763
rect 20663 22729 20697 22763
rect 21281 22729 21315 22763
rect 24777 22729 24811 22763
rect 4169 22661 4203 22695
rect 4369 22661 4403 22695
rect 7297 22661 7331 22695
rect 8769 22661 8803 22695
rect 12173 22661 12207 22695
rect 13820 22661 13854 22695
rect 17141 22661 17175 22695
rect 17258 22661 17292 22695
rect 18429 22661 18463 22695
rect 19717 22661 19751 22695
rect 20177 22661 20211 22695
rect 20453 22661 20487 22695
rect 19947 22627 19981 22661
rect 2672 22593 2706 22627
rect 3617 22593 3651 22627
rect 4896 22593 4930 22627
rect 6561 22593 6595 22627
rect 7389 22593 7423 22627
rect 8493 22593 8527 22627
rect 8585 22593 8619 22627
rect 11345 22593 11379 22627
rect 11897 22593 11931 22627
rect 11989 22593 12023 22627
rect 16037 22593 16071 22627
rect 16129 22593 16163 22627
rect 16221 22593 16255 22627
rect 16405 22593 16439 22627
rect 18337 22593 18371 22627
rect 18521 22593 18555 22627
rect 18705 22593 18739 22627
rect 18981 22593 19015 22627
rect 19257 22593 19291 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 23397 22593 23431 22627
rect 23664 22593 23698 22627
rect 25421 22593 25455 22627
rect 25605 22593 25639 22627
rect 2789 22525 2823 22559
rect 3157 22525 3191 22559
rect 3249 22525 3283 22559
rect 3709 22525 3743 22559
rect 4629 22525 4663 22559
rect 6653 22525 6687 22559
rect 6929 22525 6963 22559
rect 7180 22525 7214 22559
rect 7665 22525 7699 22559
rect 11805 22525 11839 22559
rect 13553 22525 13587 22559
rect 16773 22525 16807 22559
rect 17049 22525 17083 22559
rect 24869 22525 24903 22559
rect 8769 22457 8803 22491
rect 11529 22457 11563 22491
rect 17417 22457 17451 22491
rect 17509 22457 17543 22491
rect 18797 22457 18831 22491
rect 20913 22457 20947 22491
rect 4353 22389 4387 22423
rect 4537 22389 4571 22423
rect 6009 22389 6043 22423
rect 11253 22389 11287 22423
rect 11897 22389 11931 22423
rect 12357 22389 12391 22423
rect 17877 22389 17911 22423
rect 18061 22389 18095 22423
rect 19165 22389 19199 22423
rect 19809 22389 19843 22423
rect 19993 22389 20027 22423
rect 20637 22389 20671 22423
rect 20821 22389 20855 22423
rect 21281 22389 21315 22423
rect 21465 22389 21499 22423
rect 25789 22389 25823 22423
rect 4813 22185 4847 22219
rect 17601 22185 17635 22219
rect 17969 22185 18003 22219
rect 20085 22185 20119 22219
rect 21557 22185 21591 22219
rect 22477 22185 22511 22219
rect 24409 22185 24443 22219
rect 5273 22117 5307 22151
rect 16497 22117 16531 22151
rect 17233 22117 17267 22151
rect 18429 22117 18463 22151
rect 20637 22117 20671 22151
rect 21097 22117 21131 22151
rect 22017 22117 22051 22151
rect 2513 22049 2547 22083
rect 6009 22049 6043 22083
rect 6285 22049 6319 22083
rect 7573 22049 7607 22083
rect 10425 22049 10459 22083
rect 10609 22049 10643 22083
rect 10885 22049 10919 22083
rect 16957 22049 16991 22083
rect 20361 22049 20395 22083
rect 21373 22049 21407 22083
rect 21557 22049 21591 22083
rect 22201 22049 22235 22083
rect 24961 22049 24995 22083
rect 2421 21981 2455 22015
rect 2789 21981 2823 22015
rect 4629 21981 4663 22015
rect 4813 21981 4847 22015
rect 4905 21981 4939 22015
rect 5089 21981 5123 22015
rect 5181 21981 5215 22015
rect 5641 21981 5675 22015
rect 5917 21981 5951 22015
rect 6101 21981 6135 22015
rect 6193 21981 6227 22015
rect 6377 21981 6411 22015
rect 8309 21981 8343 22015
rect 8493 21981 8527 22015
rect 10517 21981 10551 22015
rect 10701 21981 10735 22015
rect 11437 21981 11471 22015
rect 12173 21981 12207 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 12633 21981 12667 22015
rect 12817 21981 12851 22015
rect 14105 21981 14139 22015
rect 16037 21981 16071 22015
rect 16221 21981 16255 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 17693 21981 17727 22015
rect 17877 21981 17911 22015
rect 18704 21981 18738 22015
rect 18797 21981 18831 22015
rect 21465 21981 21499 22015
rect 21925 21981 21959 22015
rect 22293 21981 22327 22015
rect 24777 21981 24811 22015
rect 25237 21981 25271 22015
rect 25605 21981 25639 22015
rect 20039 21947 20073 21981
rect 2304 21913 2338 21947
rect 5549 21913 5583 21947
rect 8058 21913 8092 21947
rect 8401 21913 8435 21947
rect 12449 21913 12483 21947
rect 20269 21913 20303 21947
rect 2145 21845 2179 21879
rect 5003 21845 5037 21879
rect 5457 21845 5491 21879
rect 5825 21845 5859 21879
rect 7849 21845 7883 21879
rect 7941 21845 7975 21879
rect 8217 21845 8251 21879
rect 10241 21845 10275 21879
rect 11621 21845 11655 21879
rect 12725 21845 12759 21879
rect 14749 21845 14783 21879
rect 16129 21845 16163 21879
rect 17417 21845 17451 21879
rect 19901 21845 19935 21879
rect 20821 21845 20855 21879
rect 20913 21845 20947 21879
rect 21833 21845 21867 21879
rect 22201 21845 22235 21879
rect 24869 21845 24903 21879
rect 25421 21845 25455 21879
rect 25789 21845 25823 21879
rect 3617 21641 3651 21675
rect 7405 21641 7439 21675
rect 7573 21641 7607 21675
rect 11345 21641 11379 21675
rect 11897 21641 11931 21675
rect 13553 21641 13587 21675
rect 22477 21641 22511 21675
rect 25145 21641 25179 21675
rect 2298 21573 2332 21607
rect 7205 21573 7239 21607
rect 20361 21573 20395 21607
rect 21557 21573 21591 21607
rect 1409 21505 1443 21539
rect 3525 21505 3559 21539
rect 3709 21505 3743 21539
rect 6837 21505 6871 21539
rect 6929 21505 6963 21539
rect 7113 21505 7147 21539
rect 7665 21505 7699 21539
rect 7932 21505 7966 21539
rect 10232 21505 10266 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 11989 21505 12023 21539
rect 12081 21505 12115 21539
rect 12348 21505 12382 21539
rect 14677 21505 14711 21539
rect 14933 21505 14967 21539
rect 19809 21505 19843 21539
rect 20085 21505 20119 21539
rect 20545 21505 20579 21539
rect 20821 21505 20855 21539
rect 21373 21505 21407 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22109 21505 22143 21539
rect 22201 21505 22235 21539
rect 22569 21505 22603 21539
rect 22845 21505 22879 21539
rect 23489 21505 23523 21539
rect 23765 21505 23799 21539
rect 24032 21505 24066 21539
rect 25789 21505 25823 21539
rect 2053 21437 2087 21471
rect 9965 21437 9999 21471
rect 15577 21437 15611 21471
rect 19901 21437 19935 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 22937 21437 22971 21471
rect 7113 21369 7147 21403
rect 19993 21369 20027 21403
rect 23673 21369 23707 21403
rect 1593 21301 1627 21335
rect 3433 21301 3467 21335
rect 7389 21301 7423 21335
rect 9045 21301 9079 21335
rect 13461 21301 13495 21335
rect 15025 21301 15059 21335
rect 20269 21301 20303 21335
rect 20637 21301 20671 21335
rect 21005 21301 21039 21335
rect 21281 21301 21315 21335
rect 25237 21301 25271 21335
rect 3341 21097 3375 21131
rect 5181 21097 5215 21131
rect 11253 21097 11287 21131
rect 13369 21097 13403 21131
rect 13553 21097 13587 21131
rect 14933 21097 14967 21131
rect 20361 21097 20395 21131
rect 20729 21097 20763 21131
rect 21833 21097 21867 21131
rect 23397 21097 23431 21131
rect 24225 21097 24259 21131
rect 5549 21029 5583 21063
rect 9505 21029 9539 21063
rect 12633 21029 12667 21063
rect 20085 21029 20119 21063
rect 6101 20961 6135 20995
rect 7205 20961 7239 20995
rect 12909 20961 12943 20995
rect 13001 20961 13035 20995
rect 13093 20961 13127 20995
rect 13645 20961 13679 20995
rect 14289 20961 14323 20995
rect 14473 20961 14507 20995
rect 15117 20961 15151 20995
rect 17233 20961 17267 20995
rect 18245 20961 18279 20995
rect 20453 20961 20487 20995
rect 21189 20961 21223 20995
rect 21557 20961 21591 20995
rect 23581 20961 23615 20995
rect 24409 20961 24443 20995
rect 1869 20893 1903 20927
rect 3341 20893 3375 20927
rect 3525 20893 3559 20927
rect 4261 20893 4295 20927
rect 4904 20893 4938 20927
rect 4997 20893 5031 20927
rect 5089 20893 5123 20927
rect 5365 20893 5399 20927
rect 5825 20893 5859 20927
rect 5917 20893 5951 20927
rect 6193 20893 6227 20927
rect 6285 20893 6319 20927
rect 7021 20893 7055 20927
rect 8769 20893 8803 20927
rect 9873 20893 9907 20927
rect 10140 20893 10174 20927
rect 11345 20893 11379 20927
rect 11529 20893 11563 20927
rect 12449 20893 12483 20927
rect 12817 20895 12851 20929
rect 13268 20893 13302 20927
rect 13921 20893 13955 20927
rect 15025 20893 15059 20927
rect 15209 20893 15243 20927
rect 17049 20893 17083 20927
rect 18061 20893 18095 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 19993 20893 20027 20927
rect 20177 20893 20211 20927
rect 20361 20893 20395 20927
rect 20821 20893 20855 20927
rect 21005 20893 21039 20927
rect 21097 20893 21131 20927
rect 21373 20893 21407 20927
rect 21649 20893 21683 20927
rect 21833 20893 21867 20927
rect 22477 20893 22511 20927
rect 22845 20893 22879 20927
rect 23029 20893 23063 20927
rect 23213 20893 23247 20927
rect 23857 20893 23891 20927
rect 2136 20825 2170 20859
rect 6653 20825 6687 20859
rect 8502 20825 8536 20859
rect 8953 20825 8987 20859
rect 9229 20825 9263 20859
rect 14565 20825 14599 20859
rect 22109 20825 22143 20859
rect 22293 20825 22327 20859
rect 23121 20825 23155 20859
rect 24676 20825 24710 20859
rect 3249 20757 3283 20791
rect 4445 20757 4479 20791
rect 4629 20757 4663 20791
rect 5641 20757 5675 20791
rect 6837 20757 6871 20791
rect 7389 20757 7423 20791
rect 9137 20757 9171 20791
rect 9321 20757 9355 20791
rect 11529 20757 11563 20791
rect 11897 20757 11931 20791
rect 16681 20757 16715 20791
rect 17141 20757 17175 20791
rect 17509 20757 17543 20791
rect 18889 20757 18923 20791
rect 19533 20757 19567 20791
rect 19809 20757 19843 20791
rect 22017 20757 22051 20791
rect 23765 20757 23799 20791
rect 25789 20757 25823 20791
rect 2053 20553 2087 20587
rect 2329 20553 2363 20587
rect 13001 20553 13035 20587
rect 13369 20553 13403 20587
rect 14013 20553 14047 20587
rect 15209 20553 15243 20587
rect 15669 20553 15703 20587
rect 16681 20553 16715 20587
rect 18153 20553 18187 20587
rect 21005 20553 21039 20587
rect 21373 20553 21407 20587
rect 23857 20553 23891 20587
rect 24685 20553 24719 20587
rect 24961 20553 24995 20587
rect 2941 20485 2975 20519
rect 3157 20485 3191 20519
rect 3433 20485 3467 20519
rect 3801 20485 3835 20519
rect 5365 20485 5399 20519
rect 8677 20485 8711 20519
rect 12642 20485 12676 20519
rect 13737 20485 13771 20519
rect 13921 20485 13955 20519
rect 17816 20485 17850 20519
rect 18521 20485 18555 20519
rect 18797 20485 18831 20519
rect 22845 20485 22879 20519
rect 23489 20485 23523 20519
rect 24317 20485 24351 20519
rect 25053 20485 25087 20519
rect 1777 20417 1811 20451
rect 1961 20417 1995 20451
rect 2421 20417 2455 20451
rect 2697 20417 2731 20451
rect 3525 20417 3559 20451
rect 3617 20417 3651 20451
rect 4445 20417 4479 20451
rect 4629 20417 4663 20451
rect 4721 20417 4755 20451
rect 4813 20417 4847 20451
rect 6193 20417 6227 20451
rect 6377 20417 6411 20451
rect 9505 20417 9539 20451
rect 9597 20417 9631 20451
rect 9781 20417 9815 20451
rect 13185 20417 13219 20451
rect 13461 20417 13495 20451
rect 14197 20417 14231 20451
rect 14381 20417 14415 20451
rect 15577 20417 15611 20451
rect 18337 20417 18371 20451
rect 18429 20417 18463 20451
rect 18705 20417 18739 20451
rect 18981 20417 19015 20451
rect 19073 20417 19107 20451
rect 19257 20417 19291 20451
rect 19349 20417 19383 20451
rect 20545 20417 20579 20451
rect 20637 20417 20671 20451
rect 20913 20417 20947 20451
rect 21189 20417 21223 20451
rect 21465 20417 21499 20451
rect 21833 20417 21867 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22385 20417 22419 20451
rect 22661 20417 22695 20451
rect 22937 20417 22971 20451
rect 23029 20417 23063 20451
rect 23305 20417 23339 20451
rect 23581 20417 23615 20451
rect 23673 20417 23707 20451
rect 24777 20417 24811 20451
rect 25697 20417 25731 20451
rect 1869 20349 1903 20383
rect 2212 20349 2246 20383
rect 3249 20349 3283 20383
rect 12909 20349 12943 20383
rect 14473 20349 14507 20383
rect 15853 20349 15887 20383
rect 18061 20349 18095 20383
rect 20821 20349 20855 20383
rect 22201 20349 22235 20383
rect 24041 20349 24075 20383
rect 24225 20349 24259 20383
rect 2789 20281 2823 20315
rect 15117 20281 15151 20315
rect 22569 20281 22603 20315
rect 23213 20281 23247 20315
rect 2973 20213 3007 20247
rect 5089 20213 5123 20247
rect 9597 20213 9631 20247
rect 11529 20213 11563 20247
rect 13553 20213 13587 20247
rect 20361 20213 20395 20247
rect 2973 20009 3007 20043
rect 4261 20009 4295 20043
rect 6377 20009 6411 20043
rect 8401 20009 8435 20043
rect 14197 20009 14231 20043
rect 17049 20009 17083 20043
rect 22201 20009 22235 20043
rect 4629 19941 4663 19975
rect 20269 19941 20303 19975
rect 22109 19941 22143 19975
rect 4353 19873 4387 19907
rect 7757 19873 7791 19907
rect 8125 19873 8159 19907
rect 15577 19873 15611 19907
rect 15669 19873 15703 19907
rect 20361 19873 20395 19907
rect 20637 19873 20671 19907
rect 20821 19873 20855 19907
rect 20913 19873 20947 19907
rect 24961 19873 24995 19907
rect 2697 19805 2731 19839
rect 2973 19805 3007 19839
rect 4261 19805 4295 19839
rect 4905 19805 4939 19839
rect 5089 19805 5123 19839
rect 5181 19805 5215 19839
rect 5365 19805 5399 19839
rect 5457 19805 5491 19839
rect 5549 19805 5583 19839
rect 6101 19805 6135 19839
rect 6469 19805 6503 19839
rect 6745 19805 6779 19839
rect 8493 19805 8527 19839
rect 8677 19805 8711 19839
rect 9045 19805 9079 19839
rect 10517 19805 10551 19839
rect 11345 19805 11379 19839
rect 11713 19805 11747 19839
rect 13737 19805 13771 19839
rect 13921 19805 13955 19839
rect 15936 19805 15970 19839
rect 18889 19805 18923 19839
rect 19257 19805 19291 19839
rect 20177 19805 20211 19839
rect 20453 19805 20487 19839
rect 21005 19805 21039 19839
rect 21097 19805 21131 19839
rect 21649 19805 21683 19839
rect 21741 19805 21775 19839
rect 21925 19805 21959 19839
rect 22569 19805 22603 19839
rect 23949 19805 23983 19839
rect 25789 19805 25823 19839
rect 6561 19737 6595 19771
rect 8242 19737 8276 19771
rect 8585 19737 8619 19771
rect 15310 19737 15344 19771
rect 18644 19737 18678 19771
rect 19993 19737 20027 19771
rect 22385 19737 22419 19771
rect 24777 19737 24811 19771
rect 25237 19737 25271 19771
rect 2789 19669 2823 19703
rect 5089 19669 5123 19703
rect 5825 19669 5859 19703
rect 5917 19669 5951 19703
rect 6929 19669 6963 19703
rect 8033 19669 8067 19703
rect 13829 19669 13863 19703
rect 17509 19669 17543 19703
rect 19901 19669 19935 19703
rect 24133 19669 24167 19703
rect 24409 19669 24443 19703
rect 24869 19669 24903 19703
rect 12909 19465 12943 19499
rect 13921 19465 13955 19499
rect 14381 19465 14415 19499
rect 14841 19465 14875 19499
rect 19073 19465 19107 19499
rect 21255 19465 21289 19499
rect 22477 19465 22511 19499
rect 23765 19465 23799 19499
rect 25237 19465 25271 19499
rect 25789 19465 25823 19499
rect 9045 19397 9079 19431
rect 10977 19397 11011 19431
rect 11774 19397 11808 19431
rect 21465 19397 21499 19431
rect 24124 19397 24158 19431
rect 2237 19329 2271 19363
rect 2697 19329 2731 19363
rect 2881 19329 2915 19363
rect 3801 19329 3835 19363
rect 4445 19329 4479 19363
rect 5549 19329 5583 19363
rect 5733 19329 5767 19363
rect 6377 19329 6411 19363
rect 6470 19329 6504 19363
rect 6653 19329 6687 19363
rect 6745 19329 6779 19363
rect 6883 19329 6917 19363
rect 8401 19329 8435 19363
rect 10701 19329 10735 19363
rect 11529 19329 11563 19363
rect 14473 19329 14507 19363
rect 15209 19329 15243 19363
rect 17233 19329 17267 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 21833 19329 21867 19363
rect 22017 19329 22051 19363
rect 22109 19329 22143 19363
rect 22201 19329 22235 19363
rect 23581 19329 23615 19363
rect 23857 19329 23891 19363
rect 25513 19329 25547 19363
rect 25605 19329 25639 19363
rect 2329 19261 2363 19295
rect 3893 19261 3927 19295
rect 4537 19261 4571 19295
rect 8493 19261 8527 19295
rect 8861 19261 8895 19295
rect 10977 19261 11011 19295
rect 13277 19261 13311 19295
rect 14565 19261 14599 19295
rect 15301 19261 15335 19295
rect 15485 19261 15519 19295
rect 17969 19261 18003 19295
rect 4169 19193 4203 19227
rect 2605 19125 2639 19159
rect 4721 19125 4755 19159
rect 5549 19125 5583 19159
rect 5917 19125 5951 19159
rect 7021 19125 7055 19159
rect 8769 19125 8803 19159
rect 10793 19125 10827 19159
rect 14013 19125 14047 19159
rect 21097 19125 21131 19159
rect 21281 19125 21315 19159
rect 25329 19125 25363 19159
rect 1593 18921 1627 18955
rect 5457 18921 5491 18955
rect 11713 18921 11747 18955
rect 12265 18921 12299 18955
rect 13829 18921 13863 18955
rect 16681 18921 16715 18955
rect 21557 18921 21591 18955
rect 23673 18921 23707 18955
rect 2697 18853 2731 18887
rect 13277 18853 13311 18887
rect 2237 18785 2271 18819
rect 3040 18785 3074 18819
rect 3157 18785 3191 18819
rect 3525 18785 3559 18819
rect 5641 18785 5675 18819
rect 8401 18785 8435 18819
rect 8585 18785 8619 18819
rect 13553 18785 13587 18819
rect 15209 18785 15243 18819
rect 17141 18785 17175 18819
rect 17325 18785 17359 18819
rect 24961 18785 24995 18819
rect 1409 18717 1443 18751
rect 2145 18717 2179 18751
rect 3249 18717 3283 18751
rect 3893 18717 3927 18751
rect 4077 18717 4111 18751
rect 4721 18717 4755 18751
rect 4813 18717 4847 18751
rect 4997 18717 5031 18751
rect 5089 18717 5123 18751
rect 5353 18717 5387 18751
rect 5825 18717 5859 18751
rect 6653 18717 6687 18751
rect 7757 18717 7791 18751
rect 8033 18717 8067 18751
rect 8309 18717 8343 18751
rect 8493 18717 8527 18751
rect 10333 18717 10367 18751
rect 12817 18717 12851 18751
rect 12909 18717 12943 18751
rect 13001 18717 13035 18751
rect 13185 18717 13219 18751
rect 13461 18717 13495 18751
rect 13921 18717 13955 18751
rect 14381 18717 14415 18751
rect 15853 18717 15887 18751
rect 17785 18717 17819 18751
rect 21189 18717 21223 18751
rect 21373 18717 21407 18751
rect 21833 18717 21867 18751
rect 21925 18695 21959 18729
rect 22293 18717 22327 18751
rect 22385 18717 22419 18751
rect 22569 18717 22603 18751
rect 22661 18717 22695 18751
rect 22753 18717 22787 18751
rect 23121 18717 23155 18751
rect 23489 18717 23523 18751
rect 25789 18717 25823 18751
rect 2697 18649 2731 18683
rect 6469 18649 6503 18683
rect 10066 18649 10100 18683
rect 11529 18649 11563 18683
rect 12081 18649 12115 18683
rect 12281 18649 12315 18683
rect 15393 18649 15427 18683
rect 22201 18649 22235 18683
rect 23305 18649 23339 18683
rect 23397 18649 23431 18683
rect 24777 18649 24811 18683
rect 25237 18649 25271 18683
rect 1961 18581 1995 18615
rect 2881 18581 2915 18615
rect 3985 18581 4019 18615
rect 5273 18581 5307 18615
rect 6009 18581 6043 18615
rect 6285 18581 6319 18615
rect 7573 18581 7607 18615
rect 7941 18581 7975 18615
rect 8769 18581 8803 18615
rect 8953 18581 8987 18615
rect 11729 18581 11763 18615
rect 11897 18581 11931 18615
rect 12449 18581 12483 18615
rect 12541 18581 12575 18615
rect 14933 18581 14967 18615
rect 15301 18581 15335 18615
rect 15761 18581 15795 18615
rect 16497 18581 16531 18615
rect 17049 18581 17083 18615
rect 18429 18581 18463 18615
rect 21649 18581 21683 18615
rect 23029 18581 23063 18615
rect 24409 18581 24443 18615
rect 24869 18581 24903 18615
rect 1869 18377 1903 18411
rect 4997 18377 5031 18411
rect 5549 18377 5583 18411
rect 8309 18377 8343 18411
rect 8677 18377 8711 18411
rect 10517 18377 10551 18411
rect 12357 18377 12391 18411
rect 12909 18377 12943 18411
rect 13553 18377 13587 18411
rect 13829 18377 13863 18411
rect 14013 18377 14047 18411
rect 14473 18377 14507 18411
rect 19809 18377 19843 18411
rect 23305 18377 23339 18411
rect 25145 18377 25179 18411
rect 25421 18377 25455 18411
rect 4353 18309 4387 18343
rect 4629 18309 4663 18343
rect 4721 18309 4755 18343
rect 10308 18309 10342 18343
rect 10425 18309 10459 18343
rect 15586 18309 15620 18343
rect 18000 18309 18034 18343
rect 18337 18309 18371 18343
rect 20269 18309 20303 18343
rect 23121 18309 23155 18343
rect 24032 18309 24066 18343
rect 2982 18241 3016 18275
rect 3249 18241 3283 18275
rect 3985 18241 4019 18275
rect 4078 18241 4112 18275
rect 4445 18241 4479 18275
rect 4813 18241 4847 18275
rect 5546 18241 5580 18275
rect 5917 18241 5951 18275
rect 6009 18241 6043 18275
rect 6929 18241 6963 18275
rect 7205 18241 7239 18275
rect 7481 18241 7515 18275
rect 7665 18241 7699 18275
rect 7849 18241 7883 18275
rect 8426 18241 8460 18275
rect 9801 18241 9835 18275
rect 12449 18241 12483 18275
rect 12725 18241 12759 18275
rect 13001 18241 13035 18275
rect 13093 18241 13127 18275
rect 13277 18241 13311 18275
rect 13369 18241 13403 18275
rect 14381 18241 14415 18275
rect 15853 18241 15887 18275
rect 18245 18241 18279 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 18889 18241 18923 18275
rect 19625 18241 19659 18275
rect 20085 18241 20119 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 20453 18241 20487 18275
rect 20545 18241 20579 18275
rect 20637 18241 20671 18275
rect 20729 18241 20763 18275
rect 20913 18241 20947 18275
rect 21557 18241 21591 18275
rect 21649 18241 21683 18275
rect 21833 18241 21867 18275
rect 21925 18241 21959 18275
rect 22293 18241 22327 18275
rect 23305 18241 23339 18275
rect 23489 18241 23523 18275
rect 23765 18241 23799 18275
rect 25237 18241 25271 18275
rect 25605 18241 25639 18275
rect 6745 18173 6779 18207
rect 7941 18173 7975 18207
rect 8217 18173 8251 18207
rect 10057 18173 10091 18207
rect 10793 18173 10827 18207
rect 11897 18173 11931 18207
rect 12633 18173 12667 18207
rect 18797 18173 18831 18207
rect 19441 18173 19475 18207
rect 19993 18173 20027 18207
rect 20821 18173 20855 18207
rect 21189 18173 21223 18207
rect 7297 18105 7331 18139
rect 8585 18105 8619 18139
rect 12265 18105 12299 18139
rect 21373 18105 21407 18139
rect 5365 18037 5399 18071
rect 7757 18037 7791 18071
rect 10149 18037 10183 18071
rect 12449 18037 12483 18071
rect 14013 18037 14047 18071
rect 16865 18037 16899 18071
rect 21833 18037 21867 18071
rect 22201 18037 22235 18071
rect 25789 18037 25823 18071
rect 2973 17833 3007 17867
rect 5457 17833 5491 17867
rect 6837 17833 6871 17867
rect 7481 17833 7515 17867
rect 8677 17833 8711 17867
rect 12449 17833 12483 17867
rect 12633 17833 12667 17867
rect 13185 17833 13219 17867
rect 14105 17833 14139 17867
rect 17877 17833 17911 17867
rect 19349 17833 19383 17867
rect 19809 17833 19843 17867
rect 21557 17833 21591 17867
rect 6377 17765 6411 17799
rect 8953 17765 8987 17799
rect 12081 17765 12115 17799
rect 13093 17765 13127 17799
rect 7113 17697 7147 17731
rect 8033 17697 8067 17731
rect 8401 17697 8435 17731
rect 8518 17697 8552 17731
rect 12725 17697 12759 17731
rect 13369 17697 13403 17731
rect 16037 17697 16071 17731
rect 16129 17697 16163 17731
rect 18337 17697 18371 17731
rect 18429 17697 18463 17731
rect 19533 17697 19567 17731
rect 21189 17697 21223 17731
rect 24961 17697 24995 17731
rect 1593 17629 1627 17663
rect 5641 17629 5675 17663
rect 5825 17629 5859 17663
rect 5917 17629 5951 17663
rect 6561 17629 6595 17663
rect 6653 17629 6687 17663
rect 7021 17629 7055 17663
rect 7205 17629 7239 17663
rect 7297 17629 7331 17663
rect 7597 17629 7631 17663
rect 7757 17629 7791 17663
rect 10066 17629 10100 17663
rect 10333 17629 10367 17663
rect 11805 17629 11839 17663
rect 13921 17629 13955 17663
rect 15485 17629 15519 17663
rect 16865 17629 16899 17663
rect 19257 17629 19291 17663
rect 19717 17629 19751 17663
rect 20821 17629 20855 17663
rect 21005 17629 21039 17663
rect 21097 17629 21131 17663
rect 21373 17629 21407 17663
rect 21833 17629 21867 17663
rect 21925 17629 21959 17663
rect 22293 17629 22327 17663
rect 25789 17629 25823 17663
rect 1860 17561 1894 17595
rect 4169 17561 4203 17595
rect 6837 17561 6871 17595
rect 8309 17561 8343 17595
rect 10609 17561 10643 17595
rect 11069 17561 11103 17595
rect 15240 17561 15274 17595
rect 17601 17561 17635 17595
rect 21649 17561 21683 17595
rect 24777 17561 24811 17595
rect 25237 17561 25271 17595
rect 4077 17493 4111 17527
rect 7665 17493 7699 17527
rect 12449 17493 12483 17527
rect 15577 17493 15611 17527
rect 15945 17493 15979 17527
rect 18245 17493 18279 17527
rect 19533 17493 19567 17527
rect 21925 17493 21959 17527
rect 24409 17493 24443 17527
rect 24869 17493 24903 17527
rect 4629 17289 4663 17323
rect 7297 17289 7331 17323
rect 8309 17289 8343 17323
rect 22201 17289 22235 17323
rect 25145 17289 25179 17323
rect 25421 17289 25455 17323
rect 7389 17221 7423 17255
rect 16865 17221 16899 17255
rect 18245 17221 18279 17255
rect 19165 17221 19199 17255
rect 20453 17221 20487 17255
rect 20545 17221 20579 17255
rect 22293 17221 22327 17255
rect 3157 17153 3191 17187
rect 4261 17153 4295 17187
rect 4415 17153 4449 17187
rect 6377 17153 6411 17187
rect 6929 17153 6963 17187
rect 7573 17153 7607 17187
rect 7665 17153 7699 17187
rect 8677 17153 8711 17187
rect 11796 17153 11830 17187
rect 13553 17153 13587 17187
rect 15229 17153 15263 17187
rect 15485 17153 15519 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 19073 17153 19107 17187
rect 19533 17153 19567 17187
rect 20269 17153 20303 17187
rect 20637 17153 20671 17187
rect 21189 17153 21223 17187
rect 21281 17153 21315 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 23305 17153 23339 17187
rect 23489 17153 23523 17187
rect 23765 17153 23799 17187
rect 24032 17153 24066 17187
rect 25237 17153 25271 17187
rect 25605 17153 25639 17187
rect 3249 17085 3283 17119
rect 3525 17085 3559 17119
rect 7021 17085 7055 17119
rect 8585 17085 8619 17119
rect 11529 17085 11563 17119
rect 16129 17085 16163 17119
rect 18337 17085 18371 17119
rect 18429 17085 18463 17119
rect 19257 17085 19291 17119
rect 20085 17085 20119 17119
rect 21097 17085 21131 17119
rect 21373 17085 21407 17119
rect 23029 17085 23063 17119
rect 7849 17017 7883 17051
rect 13001 17017 13035 17051
rect 15577 17017 15611 17051
rect 17877 17017 17911 17051
rect 25789 17017 25823 17051
rect 6469 16949 6503 16983
rect 7665 16949 7699 16983
rect 12909 16949 12943 16983
rect 14105 16949 14139 16983
rect 18705 16949 18739 16983
rect 20821 16949 20855 16983
rect 20913 16949 20947 16983
rect 22017 16949 22051 16983
rect 23673 16949 23707 16983
rect 11805 16745 11839 16779
rect 16221 16745 16255 16779
rect 18337 16745 18371 16779
rect 19901 16745 19935 16779
rect 6653 16677 6687 16711
rect 12265 16609 12299 16643
rect 12357 16609 12391 16643
rect 13461 16609 13495 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 16957 16609 16991 16643
rect 19257 16609 19291 16643
rect 20269 16609 20303 16643
rect 23581 16609 23615 16643
rect 6193 16541 6227 16575
rect 6377 16541 6411 16575
rect 17224 16541 17258 16575
rect 19993 16541 20027 16575
rect 20085 16541 20119 16575
rect 20361 16541 20395 16575
rect 20545 16541 20579 16575
rect 20821 16541 20855 16575
rect 21465 16541 21499 16575
rect 21741 16541 21775 16575
rect 21833 16541 21867 16575
rect 22109 16541 22143 16575
rect 24409 16541 24443 16575
rect 12173 16473 12207 16507
rect 20269 16473 20303 16507
rect 21925 16473 21959 16507
rect 22293 16473 22327 16507
rect 24654 16473 24688 16507
rect 12909 16405 12943 16439
rect 15853 16405 15887 16439
rect 20545 16405 20579 16439
rect 21557 16405 21591 16439
rect 23765 16405 23799 16439
rect 23857 16405 23891 16439
rect 24225 16405 24259 16439
rect 25789 16405 25823 16439
rect 1593 16201 1627 16235
rect 4445 16201 4479 16235
rect 6101 16201 6135 16235
rect 12909 16201 12943 16235
rect 18337 16201 18371 16235
rect 22845 16201 22879 16235
rect 24869 16201 24903 16235
rect 5641 16133 5675 16167
rect 6561 16133 6595 16167
rect 17224 16133 17258 16167
rect 22477 16133 22511 16167
rect 23121 16133 23155 16167
rect 1409 16065 1443 16099
rect 2329 16065 2363 16099
rect 2585 16065 2619 16099
rect 3985 16065 4019 16099
rect 4504 16065 4538 16099
rect 6377 16065 6411 16099
rect 11796 16065 11830 16099
rect 13369 16065 13403 16099
rect 13461 16065 13495 16099
rect 13829 16065 13863 16099
rect 14381 16065 14415 16099
rect 16957 16065 16991 16099
rect 19726 16065 19760 16099
rect 19993 16065 20027 16099
rect 21393 16065 21427 16099
rect 21833 16065 21867 16099
rect 22017 16065 22051 16099
rect 22293 16065 22327 16099
rect 22569 16065 22603 16099
rect 22661 16065 22695 16099
rect 22937 16065 22971 16099
rect 23213 16065 23247 16099
rect 23305 16065 23339 16099
rect 23581 16065 23615 16099
rect 23765 16065 23799 16099
rect 23857 16065 23891 16099
rect 23949 16065 23983 16099
rect 24593 16065 24627 16099
rect 25513 16065 25547 16099
rect 25605 16065 25639 16099
rect 11529 15997 11563 16031
rect 13645 15997 13679 16031
rect 21649 15997 21683 16031
rect 21925 15997 21959 16031
rect 5917 15929 5951 15963
rect 13001 15929 13035 15963
rect 24133 15929 24167 15963
rect 24777 15929 24811 15963
rect 3709 15861 3743 15895
rect 4077 15861 4111 15895
rect 4629 15861 4663 15895
rect 6745 15861 6779 15895
rect 18613 15861 18647 15895
rect 20269 15861 20303 15895
rect 23489 15861 23523 15895
rect 25789 15861 25823 15895
rect 1593 15657 1627 15691
rect 2421 15657 2455 15691
rect 2605 15657 2639 15691
rect 6929 15657 6963 15691
rect 10977 15657 11011 15691
rect 12449 15657 12483 15691
rect 18245 15657 18279 15691
rect 20177 15657 20211 15691
rect 22293 15657 22327 15691
rect 25789 15657 25823 15691
rect 17417 15589 17451 15623
rect 20637 15589 20671 15623
rect 22477 15589 22511 15623
rect 24225 15589 24259 15623
rect 12909 15521 12943 15555
rect 13093 15521 13127 15555
rect 15025 15521 15059 15555
rect 15393 15521 15427 15555
rect 17877 15521 17911 15555
rect 17969 15521 18003 15555
rect 18797 15521 18831 15555
rect 21649 15521 21683 15555
rect 22845 15521 22879 15555
rect 24961 15521 24995 15555
rect 2145 15453 2179 15487
rect 2329 15453 2363 15487
rect 2881 15453 2915 15487
rect 3065 15453 3099 15487
rect 4077 15453 4111 15487
rect 5640 15453 5674 15487
rect 5733 15453 5767 15487
rect 6561 15453 6595 15487
rect 6745 15453 6779 15487
rect 9505 15453 9539 15487
rect 10057 15453 10091 15487
rect 10241 15453 10275 15487
rect 12101 15453 12135 15487
rect 12357 15453 12391 15487
rect 14933 15453 14967 15487
rect 18705 15453 18739 15487
rect 19349 15453 19383 15487
rect 19993 15453 20027 15487
rect 20085 15453 20119 15487
rect 20545 15453 20579 15487
rect 20729 15453 20763 15487
rect 21925 15453 21959 15487
rect 22661 15453 22695 15487
rect 25237 15453 25271 15487
rect 25605 15453 25639 15487
rect 1501 15385 1535 15419
rect 2237 15385 2271 15419
rect 2573 15385 2607 15419
rect 2789 15385 2823 15419
rect 3341 15385 3375 15419
rect 3525 15385 3559 15419
rect 3985 15385 4019 15419
rect 4353 15385 4387 15419
rect 9321 15385 9355 15419
rect 9873 15385 9907 15419
rect 12817 15385 12851 15419
rect 13645 15385 13679 15419
rect 17785 15385 17819 15419
rect 23112 15385 23146 15419
rect 2973 15317 3007 15351
rect 3157 15317 3191 15351
rect 3801 15317 3835 15351
rect 4169 15317 4203 15351
rect 5365 15317 5399 15351
rect 6469 15317 6503 15351
rect 9781 15317 9815 15351
rect 10241 15317 10275 15351
rect 13369 15317 13403 15351
rect 14473 15317 14507 15351
rect 14841 15317 14875 15351
rect 15945 15317 15979 15351
rect 18613 15317 18647 15351
rect 21833 15317 21867 15351
rect 24409 15317 24443 15351
rect 25421 15317 25455 15351
rect 2789 15113 2823 15147
rect 4445 15113 4479 15147
rect 12265 15113 12299 15147
rect 15577 15113 15611 15147
rect 23305 15113 23339 15147
rect 23673 15113 23707 15147
rect 25145 15113 25179 15147
rect 1961 15045 1995 15079
rect 2973 15045 3007 15079
rect 3310 15045 3344 15079
rect 5089 15045 5123 15079
rect 5457 15045 5491 15079
rect 6377 15045 6411 15079
rect 15669 15045 15703 15079
rect 22109 15045 22143 15079
rect 23765 15045 23799 15079
rect 2605 14977 2639 15011
rect 2697 14977 2731 15011
rect 4537 14977 4571 15011
rect 4997 14977 5031 15011
rect 5181 14977 5215 15011
rect 5273 14977 5307 15011
rect 5549 14977 5583 15011
rect 5641 14977 5675 15011
rect 6745 14977 6779 15011
rect 9606 14977 9640 15011
rect 9873 14977 9907 15011
rect 9965 14977 9999 15011
rect 10232 14977 10266 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 12173 14977 12207 15011
rect 13378 14977 13412 15011
rect 13645 14977 13679 15011
rect 13737 14977 13771 15011
rect 14004 14977 14038 15011
rect 17049 14977 17083 15011
rect 17509 14977 17543 15011
rect 18061 14977 18095 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 24961 14977 24995 15011
rect 3065 14909 3099 14943
rect 6561 14909 6595 14943
rect 15761 14909 15795 14943
rect 17141 14909 17175 14943
rect 17233 14909 17267 14943
rect 23857 14909 23891 14943
rect 2329 14841 2363 14875
rect 2421 14841 2455 14875
rect 6653 14841 6687 14875
rect 8493 14841 8527 14875
rect 1777 14773 1811 14807
rect 1961 14773 1995 14807
rect 4629 14773 4663 14807
rect 5825 14773 5859 14807
rect 6561 14773 6595 14807
rect 11345 14773 11379 14807
rect 15117 14773 15151 14807
rect 15209 14773 15243 14807
rect 16681 14773 16715 14807
rect 3157 14569 3191 14603
rect 3249 14569 3283 14603
rect 4445 14569 4479 14603
rect 5641 14569 5675 14603
rect 8585 14569 8619 14603
rect 11529 14569 11563 14603
rect 11713 14569 11747 14603
rect 18797 14569 18831 14603
rect 4629 14501 4663 14535
rect 6009 14501 6043 14535
rect 8769 14501 8803 14535
rect 17141 14501 17175 14535
rect 3893 14433 3927 14467
rect 6101 14433 6135 14467
rect 13001 14433 13035 14467
rect 13921 14433 13955 14467
rect 19809 14433 19843 14467
rect 21465 14433 21499 14467
rect 1777 14365 1811 14399
rect 3433 14365 3467 14399
rect 3617 14365 3651 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4445 14365 4479 14399
rect 4721 14365 4755 14399
rect 4905 14365 4939 14399
rect 4997 14365 5031 14399
rect 5089 14365 5123 14399
rect 6285 14365 6319 14399
rect 6377 14365 6411 14399
rect 7113 14365 7147 14399
rect 7389 14365 7423 14399
rect 8953 14365 8987 14399
rect 11897 14365 11931 14399
rect 12541 14365 12575 14399
rect 12725 14365 12759 14399
rect 15402 14365 15436 14399
rect 15669 14365 15703 14399
rect 15761 14365 15795 14399
rect 17417 14365 17451 14399
rect 20545 14365 20579 14399
rect 20729 14365 20763 14399
rect 20913 14365 20947 14399
rect 21005 14365 21039 14399
rect 21097 14365 21131 14399
rect 21649 14365 21683 14399
rect 24409 14365 24443 14399
rect 2044 14297 2078 14331
rect 5365 14297 5399 14331
rect 7573 14297 7607 14331
rect 8401 14297 8435 14331
rect 9198 14297 9232 14331
rect 11345 14297 11379 14331
rect 16028 14297 16062 14331
rect 17684 14297 17718 14331
rect 21833 14297 21867 14331
rect 24654 14297 24688 14331
rect 5457 14229 5491 14263
rect 5641 14229 5675 14263
rect 6377 14229 6411 14263
rect 7205 14229 7239 14263
rect 8611 14229 8645 14263
rect 10333 14229 10367 14263
rect 11555 14229 11589 14263
rect 13277 14229 13311 14263
rect 14289 14229 14323 14263
rect 19257 14229 19291 14263
rect 19993 14229 20027 14263
rect 21373 14229 21407 14263
rect 25789 14229 25823 14263
rect 14749 14025 14783 14059
rect 16497 14025 16531 14059
rect 18521 14025 18555 14059
rect 18613 14025 18647 14059
rect 18981 14025 19015 14059
rect 19441 14025 19475 14059
rect 19809 14025 19843 14059
rect 23213 14025 23247 14059
rect 24317 14025 24351 14059
rect 25421 14025 25455 14059
rect 25789 14025 25823 14059
rect 3157 13957 3191 13991
rect 5733 13957 5767 13991
rect 6377 13957 6411 13991
rect 6577 13957 6611 13991
rect 8033 13957 8067 13991
rect 9413 13957 9447 13991
rect 9613 13957 9647 13991
rect 9965 13957 9999 13991
rect 12173 13957 12207 13991
rect 12449 13957 12483 13991
rect 12665 13957 12699 13991
rect 13001 13957 13035 13991
rect 13277 13957 13311 13991
rect 15362 13957 15396 13991
rect 17408 13957 17442 13991
rect 22078 13957 22112 13991
rect 24593 13957 24627 13991
rect 1593 13889 1627 13923
rect 1860 13889 1894 13923
rect 3065 13889 3099 13923
rect 3249 13889 3283 13923
rect 3341 13889 3375 13923
rect 3525 13889 3559 13923
rect 4905 13889 4939 13923
rect 5181 13889 5215 13923
rect 5365 13889 5399 13923
rect 5457 13889 5491 13923
rect 5549 13889 5583 13923
rect 5825 13889 5859 13923
rect 5917 13889 5951 13923
rect 7113 13889 7147 13923
rect 7389 13889 7423 13923
rect 7665 13889 7699 13923
rect 7757 13889 7791 13923
rect 8308 13911 8342 13945
rect 8401 13887 8435 13921
rect 8585 13889 8619 13923
rect 8683 13889 8717 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 9045 13889 9079 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 11805 13889 11839 13923
rect 13093 13889 13127 13923
rect 15117 13889 15151 13923
rect 17141 13889 17175 13923
rect 19073 13889 19107 13923
rect 19901 13889 19935 13923
rect 20269 13889 20303 13923
rect 20525 13889 20559 13923
rect 21833 13889 21867 13923
rect 23673 13889 23707 13923
rect 23857 13889 23891 13923
rect 23949 13889 23983 13923
rect 24041 13889 24075 13923
rect 24409 13889 24443 13923
rect 25237 13889 25271 13923
rect 25605 13889 25639 13923
rect 5273 13821 5307 13855
rect 8033 13821 8067 13855
rect 19165 13821 19199 13855
rect 19993 13821 20027 13855
rect 24777 13821 24811 13855
rect 2973 13753 3007 13787
rect 6101 13753 6135 13787
rect 6745 13753 6779 13787
rect 7297 13753 7331 13787
rect 9781 13753 9815 13787
rect 12357 13753 12391 13787
rect 12817 13753 12851 13787
rect 21649 13753 21683 13787
rect 3341 13685 3375 13719
rect 4997 13685 5031 13719
rect 6561 13685 6595 13719
rect 8217 13685 8251 13719
rect 8493 13685 8527 13719
rect 9321 13685 9355 13719
rect 9597 13685 9631 13719
rect 12173 13685 12207 13719
rect 12633 13685 12667 13719
rect 2145 13481 2179 13515
rect 2329 13481 2363 13515
rect 5181 13481 5215 13515
rect 6285 13481 6319 13515
rect 7113 13481 7147 13515
rect 7481 13481 7515 13515
rect 8217 13481 8251 13515
rect 8677 13481 8711 13515
rect 9229 13481 9263 13515
rect 13921 13481 13955 13515
rect 15577 13481 15611 13515
rect 18521 13481 18555 13515
rect 20177 13481 20211 13515
rect 5457 13413 5491 13447
rect 5549 13413 5583 13447
rect 6929 13413 6963 13447
rect 7640 13345 7674 13379
rect 13369 13345 13403 13379
rect 14933 13345 14967 13379
rect 16221 13345 16255 13379
rect 17141 13345 17175 13379
rect 19809 13345 19843 13379
rect 20913 13345 20947 13379
rect 23489 13345 23523 13379
rect 5365 13277 5399 13311
rect 5641 13277 5675 13311
rect 5825 13277 5859 13311
rect 5917 13277 5951 13311
rect 6101 13277 6135 13311
rect 7113 13277 7147 13311
rect 7205 13277 7239 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 8493 13277 8527 13311
rect 8769 13277 8803 13311
rect 8953 13277 8987 13311
rect 12265 13277 12299 13311
rect 12449 13277 12483 13311
rect 13553 13277 13587 13311
rect 20453 13277 20487 13311
rect 20545 13277 20579 13311
rect 20637 13277 20671 13311
rect 20821 13277 20855 13311
rect 23581 13277 23615 13311
rect 23765 13277 23799 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 24409 13277 24443 13311
rect 2513 13209 2547 13243
rect 7389 13209 7423 13243
rect 9229 13209 9263 13243
rect 13461 13209 13495 13243
rect 15117 13209 15151 13243
rect 17408 13209 17442 13243
rect 21180 13209 21214 13243
rect 22385 13209 22419 13243
rect 22569 13209 22603 13243
rect 23121 13209 23155 13243
rect 23305 13209 23339 13243
rect 24225 13209 24259 13243
rect 24654 13209 24688 13243
rect 2313 13141 2347 13175
rect 9045 13141 9079 13175
rect 12081 13141 12115 13175
rect 15209 13141 15243 13175
rect 15669 13141 15703 13175
rect 19257 13141 19291 13175
rect 22293 13141 22327 13175
rect 22753 13141 22787 13175
rect 25789 13141 25823 13175
rect 5089 12937 5123 12971
rect 8033 12937 8067 12971
rect 8125 12937 8159 12971
rect 9137 12937 9171 12971
rect 17877 12937 17911 12971
rect 18245 12937 18279 12971
rect 19533 12937 19567 12971
rect 21189 12937 21223 12971
rect 21281 12937 21315 12971
rect 25789 12937 25823 12971
rect 5549 12869 5583 12903
rect 7665 12869 7699 12903
rect 8309 12869 8343 12903
rect 8769 12869 8803 12903
rect 8969 12869 9003 12903
rect 10342 12869 10376 12903
rect 23765 12869 23799 12903
rect 2881 12801 2915 12835
rect 3065 12801 3099 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 7849 12801 7883 12835
rect 8493 12801 8527 12835
rect 11980 12801 12014 12835
rect 18337 12801 18371 12835
rect 19717 12801 19751 12835
rect 19809 12801 19843 12835
rect 19993 12801 20027 12835
rect 20085 12801 20119 12835
rect 20545 12801 20579 12835
rect 20729 12801 20763 12835
rect 20821 12801 20855 12835
rect 20913 12801 20947 12835
rect 21465 12801 21499 12835
rect 21649 12801 21683 12835
rect 23581 12801 23615 12835
rect 23673 12801 23707 12835
rect 23949 12801 23983 12835
rect 24041 12801 24075 12835
rect 24308 12801 24342 12835
rect 25611 12801 25645 12835
rect 5089 12733 5123 12767
rect 10609 12733 10643 12767
rect 11713 12733 11747 12767
rect 18429 12733 18463 12767
rect 5733 12665 5767 12699
rect 3065 12597 3099 12631
rect 5273 12597 5307 12631
rect 8953 12597 8987 12631
rect 9229 12597 9263 12631
rect 13093 12597 13127 12631
rect 23397 12597 23431 12631
rect 25421 12597 25455 12631
rect 3433 12393 3467 12427
rect 5181 12393 5215 12427
rect 8953 12393 8987 12427
rect 19901 12393 19935 12427
rect 20545 12393 20579 12427
rect 25053 12393 25087 12427
rect 25145 12393 25179 12427
rect 12909 12325 12943 12359
rect 22017 12325 22051 12359
rect 9229 12257 9263 12291
rect 11345 12257 11379 12291
rect 13461 12257 13495 12291
rect 16221 12257 16255 12291
rect 17877 12257 17911 12291
rect 2329 12189 2363 12223
rect 2789 12189 2823 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 5457 12189 5491 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 8769 12189 8803 12223
rect 9321 12189 9355 12223
rect 11612 12189 11646 12223
rect 13277 12189 13311 12223
rect 14105 12189 14139 12223
rect 18797 12189 18831 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 20361 12189 20395 12223
rect 20453 12189 20487 12223
rect 20729 12189 20763 12223
rect 20821 12189 20855 12223
rect 21005 12189 21039 12223
rect 21097 12189 21131 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 22201 12189 22235 12223
rect 22385 12189 22419 12223
rect 22569 12189 22603 12223
rect 24409 12189 24443 12223
rect 24593 12189 24627 12223
rect 24685 12189 24719 12223
rect 24777 12189 24811 12223
rect 25329 12189 25363 12223
rect 25513 12189 25547 12223
rect 25697 12189 25731 12223
rect 2697 12121 2731 12155
rect 2973 12121 3007 12155
rect 3157 12121 3191 12155
rect 3412 12121 3446 12155
rect 3617 12121 3651 12155
rect 5181 12121 5215 12155
rect 8401 12121 8435 12155
rect 14372 12121 14406 12155
rect 17693 12121 17727 12155
rect 18153 12121 18187 12155
rect 22293 12121 22327 12155
rect 23857 12121 23891 12155
rect 24041 12121 24075 12155
rect 24225 12121 24259 12155
rect 25421 12121 25455 12155
rect 2145 12053 2179 12087
rect 2421 12053 2455 12087
rect 2513 12053 2547 12087
rect 3249 12053 3283 12087
rect 3893 12053 3927 12087
rect 5365 12053 5399 12087
rect 8677 12053 8711 12087
rect 12725 12053 12759 12087
rect 13369 12053 13403 12087
rect 15485 12053 15519 12087
rect 15669 12053 15703 12087
rect 16037 12053 16071 12087
rect 16129 12053 16163 12087
rect 17325 12053 17359 12087
rect 17785 12053 17819 12087
rect 21189 12053 21223 12087
rect 1593 11849 1627 11883
rect 3157 11849 3191 11883
rect 3325 11849 3359 11883
rect 4353 11849 4387 11883
rect 5089 11849 5123 11883
rect 5733 11849 5767 11883
rect 7849 11849 7883 11883
rect 8309 11849 8343 11883
rect 12909 11849 12943 11883
rect 13093 11849 13127 11883
rect 14657 11849 14691 11883
rect 18429 11849 18463 11883
rect 21005 11849 21039 11883
rect 25789 11849 25823 11883
rect 3525 11781 3559 11815
rect 3893 11781 3927 11815
rect 8217 11781 8251 11815
rect 13645 11781 13679 11815
rect 17316 11781 17350 11815
rect 1409 11713 1443 11747
rect 1593 11713 1627 11747
rect 1685 11713 1719 11747
rect 1952 11713 1986 11747
rect 3801 11713 3835 11747
rect 3985 11713 4019 11747
rect 4261 11713 4295 11747
rect 4537 11713 4571 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 5181 11713 5215 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 7941 11713 7975 11747
rect 8033 11713 8067 11747
rect 9422 11713 9456 11747
rect 9689 11713 9723 11747
rect 11529 11713 11563 11747
rect 11796 11713 11830 11747
rect 13001 11713 13035 11747
rect 13185 11713 13219 11747
rect 13277 11713 13311 11747
rect 14289 11713 14323 11747
rect 14749 11713 14783 11747
rect 15016 11713 15050 11747
rect 17049 11713 17083 11747
rect 18889 11713 18923 11747
rect 19625 11713 19659 11747
rect 19892 11713 19926 11747
rect 21189 11713 21223 11747
rect 21833 11713 21867 11747
rect 22089 11713 22123 11747
rect 24124 11713 24158 11747
rect 25605 11713 25639 11747
rect 4629 11645 4663 11679
rect 7665 11645 7699 11679
rect 14013 11645 14047 11679
rect 14197 11645 14231 11679
rect 18981 11645 19015 11679
rect 19073 11645 19107 11679
rect 23857 11645 23891 11679
rect 3617 11577 3651 11611
rect 4169 11577 4203 11611
rect 5273 11577 5307 11611
rect 13829 11577 13863 11611
rect 25237 11577 25271 11611
rect 3065 11509 3099 11543
rect 3341 11509 3375 11543
rect 4537 11509 4571 11543
rect 13645 11509 13679 11543
rect 16129 11509 16163 11543
rect 18521 11509 18555 11543
rect 21281 11509 21315 11543
rect 23213 11509 23247 11543
rect 3433 11305 3467 11339
rect 3985 11305 4019 11339
rect 5273 11305 5307 11339
rect 6745 11305 6779 11339
rect 7389 11305 7423 11339
rect 7849 11305 7883 11339
rect 8033 11305 8067 11339
rect 8585 11305 8619 11339
rect 8769 11305 8803 11339
rect 11989 11305 12023 11339
rect 12909 11305 12943 11339
rect 14289 11305 14323 11339
rect 14749 11305 14783 11339
rect 15016 11305 15050 11339
rect 18705 11305 18739 11339
rect 19257 11305 19291 11339
rect 19993 11305 20027 11339
rect 21741 11305 21775 11339
rect 25789 11305 25823 11339
rect 7113 11237 7147 11271
rect 7573 11237 7607 11271
rect 20729 11237 20763 11271
rect 24869 11237 24903 11271
rect 4353 11169 4387 11203
rect 4997 11169 5031 11203
rect 14473 11169 14507 11203
rect 15301 11169 15335 11203
rect 17325 11169 17359 11203
rect 19809 11169 19843 11203
rect 22477 11169 22511 11203
rect 24225 11169 24259 11203
rect 2053 11101 2087 11135
rect 4261 11101 4295 11135
rect 4445 11101 4479 11135
rect 4905 11101 4939 11135
rect 5365 11101 5399 11135
rect 6837 11101 6871 11135
rect 8125 11101 8159 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 12173 11101 12207 11135
rect 12633 11101 12667 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 14197 11101 14231 11135
rect 17592 11101 17626 11135
rect 20269 11101 20303 11135
rect 20361 11101 20395 11135
rect 20453 11101 20487 11135
rect 20637 11101 20671 11135
rect 20913 11101 20947 11135
rect 21005 11101 21039 11135
rect 21189 11101 21223 11135
rect 21281 11101 21315 11135
rect 22017 11101 22051 11135
rect 22109 11101 22143 11135
rect 22201 11101 22235 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 23581 11101 23615 11135
rect 23765 11101 23799 11135
rect 23857 11101 23891 11135
rect 23949 11101 23983 11135
rect 24777 11101 24811 11135
rect 25605 11101 25639 11135
rect 2320 11033 2354 11067
rect 3801 11033 3835 11067
rect 4006 11033 4040 11067
rect 5632 11033 5666 11067
rect 6929 11033 6963 11067
rect 7113 11033 7147 11067
rect 7205 11033 7239 11067
rect 7405 11033 7439 11067
rect 7665 11033 7699 11067
rect 8401 11033 8435 11067
rect 8617 11033 8651 11067
rect 12357 11033 12391 11067
rect 12449 11033 12483 11067
rect 14841 11033 14875 11067
rect 15546 11033 15580 11067
rect 22845 11033 22879 11067
rect 24409 11033 24443 11067
rect 24593 11033 24627 11067
rect 25053 11033 25087 11067
rect 25237 11033 25271 11067
rect 4169 10965 4203 10999
rect 7875 10965 7909 10999
rect 15041 10965 15075 10999
rect 15209 10965 15243 10999
rect 16681 10965 16715 10999
rect 2881 10761 2915 10795
rect 5457 10761 5491 10795
rect 7205 10761 7239 10795
rect 7573 10761 7607 10795
rect 11621 10761 11655 10795
rect 12633 10761 12667 10795
rect 14381 10761 14415 10795
rect 15393 10761 15427 10795
rect 25789 10761 25823 10795
rect 5609 10693 5643 10727
rect 5825 10693 5859 10727
rect 8686 10693 8720 10727
rect 10977 10693 11011 10727
rect 21833 10693 21867 10727
rect 22017 10693 22051 10727
rect 22201 10693 22235 10727
rect 24041 10693 24075 10727
rect 24378 10693 24412 10727
rect 4005 10625 4039 10659
rect 4261 10625 4295 10659
rect 6837 10625 6871 10659
rect 8953 10625 8987 10659
rect 10241 10625 10275 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 12081 10625 12115 10659
rect 12265 10625 12299 10659
rect 12449 10625 12483 10659
rect 12633 10625 12667 10659
rect 14289 10625 14323 10659
rect 14565 10625 14599 10659
rect 14841 10625 14875 10659
rect 15761 10625 15795 10659
rect 18337 10625 18371 10659
rect 21281 10625 21315 10659
rect 21373 10625 21407 10659
rect 21465 10625 21499 10659
rect 21649 10625 21683 10659
rect 23397 10625 23431 10659
rect 23581 10625 23615 10659
rect 23673 10625 23707 10659
rect 23765 10625 23799 10659
rect 25605 10625 25639 10659
rect 6745 10557 6779 10591
rect 15853 10557 15887 10591
rect 15945 10557 15979 10591
rect 18429 10557 18463 10591
rect 18613 10557 18647 10591
rect 24133 10557 24167 10591
rect 5641 10421 5675 10455
rect 12173 10421 12207 10455
rect 14657 10421 14691 10455
rect 15117 10421 15151 10455
rect 17969 10421 18003 10455
rect 21005 10421 21039 10455
rect 25513 10421 25547 10455
rect 12725 10217 12759 10251
rect 13645 10217 13679 10251
rect 14197 10217 14231 10251
rect 14749 10217 14783 10251
rect 18981 10217 19015 10251
rect 24409 10217 24443 10251
rect 25789 10217 25823 10251
rect 15209 10149 15243 10183
rect 22293 10149 22327 10183
rect 15945 10081 15979 10115
rect 19809 10081 19843 10115
rect 20913 10081 20947 10115
rect 3617 10013 3651 10047
rect 3893 10013 3927 10047
rect 4721 10013 4755 10047
rect 9689 10013 9723 10047
rect 9873 10013 9907 10047
rect 10425 10013 10459 10047
rect 13369 10013 13403 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14657 10013 14691 10047
rect 14933 10013 14967 10047
rect 17601 10013 17635 10047
rect 17868 10013 17902 10047
rect 20637 10013 20671 10047
rect 21169 10013 21203 10047
rect 24593 10013 24627 10047
rect 24685 10013 24719 10047
rect 24961 10013 24995 10047
rect 25237 10013 25271 10047
rect 25605 10013 25639 10047
rect 13613 9945 13647 9979
rect 13829 9945 13863 9979
rect 15761 9945 15795 9979
rect 19625 9945 19659 9979
rect 20085 9945 20119 9979
rect 24777 9945 24811 9979
rect 9781 9877 9815 9911
rect 13461 9877 13495 9911
rect 14473 9877 14507 9911
rect 15393 9877 15427 9911
rect 15853 9877 15887 9911
rect 19257 9877 19291 9911
rect 19717 9877 19751 9911
rect 25421 9877 25455 9911
rect 19625 9673 19659 9707
rect 22109 9673 22143 9707
rect 3309 9605 3343 9639
rect 3525 9605 3559 9639
rect 11796 9605 11830 9639
rect 14473 9605 14507 9639
rect 15292 9605 15326 9639
rect 17868 9605 17902 9639
rect 23765 9605 23799 9639
rect 24102 9605 24136 9639
rect 4077 9537 4111 9571
rect 9965 9537 9999 9571
rect 10232 9537 10266 9571
rect 11529 9537 11563 9571
rect 15025 9537 15059 9571
rect 17049 9537 17083 9571
rect 19349 9537 19383 9571
rect 19717 9537 19751 9571
rect 21925 9537 21959 9571
rect 23121 9537 23155 9571
rect 23305 9537 23339 9571
rect 23397 9537 23431 9571
rect 23489 9537 23523 9571
rect 23857 9537 23891 9571
rect 9321 9469 9355 9503
rect 13001 9469 13035 9503
rect 14565 9469 14599 9503
rect 14657 9469 14691 9503
rect 17141 9469 17175 9503
rect 17233 9469 17267 9503
rect 17601 9469 17635 9503
rect 19257 9469 19291 9503
rect 16405 9401 16439 9435
rect 18981 9401 19015 9435
rect 3157 9333 3191 9367
rect 3341 9333 3375 9367
rect 9873 9333 9907 9367
rect 11345 9333 11379 9367
rect 12909 9333 12943 9367
rect 13645 9333 13679 9367
rect 14105 9333 14139 9367
rect 16681 9333 16715 9367
rect 25237 9333 25271 9367
rect 1685 9129 1719 9163
rect 13277 9129 13311 9163
rect 13645 9129 13679 9163
rect 16589 9129 16623 9163
rect 19441 9129 19475 9163
rect 22569 9129 22603 9163
rect 24777 9129 24811 9163
rect 6009 9061 6043 9095
rect 6653 9061 6687 9095
rect 7205 9061 7239 9095
rect 9229 9061 9263 9095
rect 22477 9061 22511 9095
rect 6745 8993 6779 9027
rect 12173 8993 12207 9027
rect 12290 8993 12324 9027
rect 13185 8993 13219 9027
rect 15209 8993 15243 9027
rect 21097 8993 21131 9027
rect 2798 8925 2832 8959
rect 3065 8925 3099 8959
rect 3157 8925 3191 8959
rect 3433 8925 3467 8959
rect 4077 8925 4111 8959
rect 5273 8925 5307 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 5733 8925 5767 8959
rect 6469 8925 6503 8959
rect 6837 8925 6871 8959
rect 6930 8925 6964 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 11805 8925 11839 8959
rect 13277 8925 13311 8959
rect 13461 8925 13495 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 15476 8925 15510 8959
rect 18981 8925 19015 8959
rect 20637 8925 20671 8959
rect 20729 8925 20763 8959
rect 20821 8925 20855 8959
rect 21005 8925 21039 8959
rect 22753 8925 22787 8959
rect 24409 8925 24443 8959
rect 24593 8925 24627 8959
rect 25605 8925 25639 8959
rect 4905 8857 4939 8891
rect 5089 8857 5123 8891
rect 5641 8857 5675 8891
rect 6285 8857 6319 8891
rect 9229 8857 9263 8891
rect 9566 8857 9600 8891
rect 10793 8857 10827 8891
rect 12081 8857 12115 8891
rect 14197 8857 14231 8891
rect 19257 8857 19291 8891
rect 19441 8857 19475 8891
rect 20361 8857 20395 8891
rect 21342 8857 21376 8891
rect 22937 8857 22971 8891
rect 25053 8857 25087 8891
rect 25237 8857 25271 8891
rect 3249 8789 3283 8823
rect 3617 8789 3651 8823
rect 6193 8789 6227 8823
rect 9045 8789 9079 8823
rect 10701 8789 10735 8823
rect 12449 8789 12483 8823
rect 12541 8789 12575 8823
rect 18889 8789 18923 8823
rect 19625 8789 19659 8823
rect 24869 8789 24903 8823
rect 25789 8789 25823 8823
rect 1777 8585 1811 8619
rect 2605 8585 2639 8619
rect 2789 8585 2823 8619
rect 4721 8585 4755 8619
rect 6193 8585 6227 8619
rect 11345 8585 11379 8619
rect 18521 8585 18555 8619
rect 19809 8585 19843 8619
rect 23765 8585 23799 8619
rect 1961 8517 1995 8551
rect 2145 8517 2179 8551
rect 4537 8517 4571 8551
rect 7941 8517 7975 8551
rect 8125 8517 8159 8551
rect 9689 8517 9723 8551
rect 13001 8517 13035 8551
rect 16037 8517 16071 8551
rect 17417 8517 17451 8551
rect 17785 8517 17819 8551
rect 18705 8517 18739 8551
rect 22569 8517 22603 8551
rect 24102 8517 24136 8551
rect 25697 8517 25731 8551
rect 3148 8449 3182 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 5080 8449 5114 8483
rect 6561 8449 6595 8483
rect 6929 8449 6963 8483
rect 7113 8449 7147 8483
rect 7849 8449 7883 8483
rect 8217 8449 8251 8483
rect 8473 8449 8507 8483
rect 11529 8449 11563 8483
rect 11785 8449 11819 8483
rect 13185 8449 13219 8483
rect 13369 8449 13403 8483
rect 13461 8449 13495 8483
rect 13553 8449 13587 8483
rect 13829 8449 13863 8483
rect 14096 8449 14130 8483
rect 16681 8449 16715 8483
rect 17693 8449 17727 8483
rect 19073 8449 19107 8483
rect 19625 8449 19659 8483
rect 20085 8449 20119 8483
rect 20269 8449 20303 8483
rect 21373 8449 21407 8483
rect 21557 8449 21591 8483
rect 22017 8449 22051 8483
rect 22109 8449 22143 8483
rect 22201 8449 22235 8483
rect 22385 8449 22419 8483
rect 23121 8449 23155 8483
rect 23305 8449 23339 8483
rect 23397 8449 23431 8483
rect 23489 8449 23523 8483
rect 23857 8449 23891 8483
rect 25329 8449 25363 8483
rect 25513 8449 25547 8483
rect 2237 8381 2271 8415
rect 2881 8381 2915 8415
rect 6837 8381 6871 8415
rect 10517 8381 10551 8415
rect 10793 8381 10827 8415
rect 13737 8381 13771 8415
rect 18981 8381 19015 8415
rect 8125 8313 8159 8347
rect 9597 8313 9631 8347
rect 15209 8313 15243 8347
rect 18337 8313 18371 8347
rect 21557 8313 21591 8347
rect 25237 8313 25271 8347
rect 2605 8245 2639 8279
rect 4261 8245 4295 8279
rect 6377 8245 6411 8279
rect 6745 8245 6779 8279
rect 7297 8245 7331 8279
rect 12909 8245 12943 8279
rect 13645 8245 13679 8279
rect 18521 8245 18555 8279
rect 21833 8245 21867 8279
rect 2421 8041 2455 8075
rect 3157 8041 3191 8075
rect 5641 8041 5675 8075
rect 5825 8041 5859 8075
rect 7665 8041 7699 8075
rect 11713 8041 11747 8075
rect 11989 8041 12023 8075
rect 12173 8041 12207 8075
rect 17417 8041 17451 8075
rect 19349 8041 19383 8075
rect 2973 7973 3007 8007
rect 6193 7973 6227 8007
rect 7481 7973 7515 8007
rect 8953 7973 8987 8007
rect 13921 7973 13955 8007
rect 18061 7973 18095 8007
rect 4353 7905 4387 7939
rect 5181 7905 5215 7939
rect 8033 7905 8067 7939
rect 8217 7905 8251 7939
rect 11161 7905 11195 7939
rect 13093 7905 13127 7939
rect 13369 7905 13403 7939
rect 24409 7905 24443 7939
rect 2789 7837 2823 7871
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3341 7837 3375 7871
rect 3525 7837 3559 7871
rect 3617 7837 3651 7871
rect 3893 7837 3927 7871
rect 3985 7837 4019 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 4997 7837 5031 7871
rect 5089 7837 5123 7871
rect 5365 7837 5399 7871
rect 6561 7837 6595 7871
rect 6654 7837 6688 7871
rect 6929 7837 6963 7871
rect 7067 7837 7101 7871
rect 10333 7837 10367 7871
rect 10885 7837 10919 7871
rect 11069 7837 11103 7871
rect 11805 7837 11839 7871
rect 11897 7837 11931 7871
rect 14105 7837 14139 7871
rect 17509 7837 17543 7871
rect 17877 7837 17911 7871
rect 17969 7837 18003 7871
rect 18245 7837 18279 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 19257 7837 19291 7871
rect 19533 7837 19567 7871
rect 20729 7837 20763 7871
rect 22937 7837 22971 7871
rect 23213 7837 23247 7871
rect 23397 7837 23431 7871
rect 23489 7837 23523 7871
rect 23581 7837 23615 7871
rect 2421 7769 2455 7803
rect 6837 7769 6871 7803
rect 10088 7769 10122 7803
rect 10701 7769 10735 7803
rect 12141 7769 12175 7803
rect 12357 7769 12391 7803
rect 13461 7769 13495 7803
rect 14350 7769 14384 7803
rect 16129 7769 16163 7803
rect 17693 7769 17727 7803
rect 18337 7769 18371 7803
rect 20996 7769 21030 7803
rect 22201 7769 22235 7803
rect 24654 7769 24688 7803
rect 2237 7701 2271 7735
rect 5549 7701 5583 7735
rect 5825 7701 5859 7735
rect 7205 7701 7239 7735
rect 7665 7701 7699 7735
rect 8769 7701 8803 7735
rect 11529 7701 11563 7735
rect 12449 7701 12483 7735
rect 13553 7701 13587 7735
rect 15485 7701 15519 7735
rect 19073 7701 19107 7735
rect 22109 7701 22143 7735
rect 23857 7701 23891 7735
rect 25789 7701 25823 7735
rect 3893 7497 3927 7531
rect 4353 7497 4387 7531
rect 7389 7497 7423 7531
rect 8033 7497 8067 7531
rect 9137 7497 9171 7531
rect 10701 7497 10735 7531
rect 12173 7497 12207 7531
rect 16681 7497 16715 7531
rect 20821 7497 20855 7531
rect 25329 7497 25363 7531
rect 25789 7497 25823 7531
rect 4045 7429 4079 7463
rect 4261 7429 4295 7463
rect 8953 7429 8987 7463
rect 19625 7429 19659 7463
rect 21833 7429 21867 7463
rect 24194 7429 24228 7463
rect 2320 7361 2354 7395
rect 4537 7361 4571 7395
rect 6837 7361 6871 7395
rect 7002 7361 7036 7395
rect 7113 7361 7147 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 7941 7361 7975 7395
rect 8217 7361 8251 7395
rect 8677 7361 8711 7395
rect 8769 7361 8803 7395
rect 10425 7361 10459 7395
rect 10517 7361 10551 7395
rect 10977 7361 11011 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 12725 7361 12759 7395
rect 15117 7361 15151 7395
rect 15384 7361 15418 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 17141 7361 17175 7395
rect 17233 7361 17267 7395
rect 19165 7361 19199 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 19533 7361 19567 7395
rect 19809 7361 19843 7395
rect 19993 7361 20027 7395
rect 20361 7361 20395 7395
rect 20545 7361 20579 7395
rect 21097 7361 21131 7395
rect 21189 7361 21223 7395
rect 21281 7361 21315 7395
rect 21465 7361 21499 7395
rect 23213 7361 23247 7395
rect 23397 7361 23431 7395
rect 23489 7361 23523 7395
rect 23581 7361 23615 7395
rect 23949 7361 23983 7395
rect 25605 7361 25639 7395
rect 2053 7293 2087 7327
rect 4721 7293 4755 7327
rect 8309 7293 8343 7327
rect 10701 7293 10735 7327
rect 11069 7293 11103 7327
rect 11989 7293 12023 7327
rect 12357 7293 12391 7327
rect 12449 7293 12483 7327
rect 12633 7293 12667 7327
rect 22661 7293 22695 7327
rect 23857 7293 23891 7327
rect 11345 7225 11379 7259
rect 11621 7225 11655 7259
rect 12541 7225 12575 7259
rect 3433 7157 3467 7191
rect 4077 7157 4111 7191
rect 8585 7157 8619 7191
rect 11989 7157 12023 7191
rect 16497 7157 16531 7191
rect 18889 7157 18923 7191
rect 20729 7157 20763 7191
rect 7389 6953 7423 6987
rect 10793 6953 10827 6987
rect 12449 6953 12483 6987
rect 14933 6953 14967 6987
rect 17969 6885 18003 6919
rect 1961 6817 1995 6851
rect 4353 6817 4387 6851
rect 8953 6817 8987 6851
rect 10977 6817 11011 6851
rect 22661 6817 22695 6851
rect 23489 6817 23523 6851
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 7113 6749 7147 6783
rect 8769 6749 8803 6783
rect 9597 6749 9631 6783
rect 9689 6749 9723 6783
rect 10701 6749 10735 6783
rect 11069 6749 11103 6783
rect 11336 6749 11370 6783
rect 14105 6749 14139 6783
rect 15117 6749 15151 6783
rect 15209 6749 15243 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 16681 6749 16715 6783
rect 17141 6749 17175 6783
rect 18417 6749 18451 6783
rect 18613 6749 18647 6783
rect 18705 6749 18739 6783
rect 18797 6749 18831 6783
rect 19257 6749 19291 6783
rect 20729 6749 20763 6783
rect 20913 6749 20947 6783
rect 21005 6749 21039 6783
rect 21097 6749 21131 6783
rect 22201 6749 22235 6783
rect 22385 6749 22419 6783
rect 22569 6749 22603 6783
rect 23673 6749 23707 6783
rect 24593 6749 24627 6783
rect 24685 6749 24719 6783
rect 24961 6749 24995 6783
rect 25237 6749 25271 6783
rect 25605 6749 25639 6783
rect 2228 6681 2262 6715
rect 3801 6681 3835 6715
rect 4077 6681 4111 6715
rect 8524 6681 8558 6715
rect 14289 6681 14323 6715
rect 15853 6681 15887 6715
rect 16957 6681 16991 6715
rect 18153 6681 18187 6715
rect 18337 6681 18371 6715
rect 19073 6681 19107 6715
rect 19502 6681 19536 6715
rect 22845 6681 22879 6715
rect 23029 6681 23063 6715
rect 23857 6681 23891 6715
rect 24777 6681 24811 6715
rect 3341 6613 3375 6647
rect 7205 6613 7239 6647
rect 9781 6613 9815 6647
rect 10977 6613 11011 6647
rect 14473 6613 14507 6647
rect 16773 6613 16807 6647
rect 20637 6613 20671 6647
rect 21373 6613 21407 6647
rect 24409 6613 24443 6647
rect 25421 6613 25455 6647
rect 25789 6613 25823 6647
rect 2237 6409 2271 6443
rect 2329 6409 2363 6443
rect 2789 6409 2823 6443
rect 3893 6409 3927 6443
rect 6009 6409 6043 6443
rect 8125 6409 8159 6443
rect 8953 6409 8987 6443
rect 15577 6409 15611 6443
rect 16681 6409 16715 6443
rect 2145 6341 2179 6375
rect 2481 6341 2515 6375
rect 2697 6341 2731 6375
rect 5181 6341 5215 6375
rect 5381 6341 5415 6375
rect 9045 6341 9079 6375
rect 9413 6341 9447 6375
rect 9657 6341 9691 6375
rect 9873 6341 9907 6375
rect 11069 6341 11103 6375
rect 19340 6341 19374 6375
rect 23581 6341 23615 6375
rect 23918 6341 23952 6375
rect 25421 6341 25455 6375
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 3065 6273 3099 6307
rect 3157 6273 3191 6307
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 3525 6273 3559 6307
rect 3709 6273 3743 6307
rect 5825 6273 5859 6307
rect 6101 6273 6135 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7389 6273 7423 6307
rect 7481 6273 7515 6307
rect 7757 6273 7791 6307
rect 8217 6273 8251 6307
rect 9229 6273 9263 6307
rect 10885 6273 10919 6307
rect 10977 6273 11011 6307
rect 11207 6273 11241 6307
rect 11805 6273 11839 6307
rect 13277 6273 13311 6307
rect 13544 6273 13578 6307
rect 15853 6273 15887 6307
rect 15945 6273 15979 6307
rect 16037 6273 16071 6307
rect 16221 6273 16255 6307
rect 16865 6273 16899 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 17233 6273 17267 6307
rect 21281 6273 21315 6307
rect 21373 6273 21407 6307
rect 22937 6273 22971 6307
rect 23121 6273 23155 6307
rect 23213 6273 23247 6307
rect 23305 6273 23339 6307
rect 25329 6273 25363 6307
rect 25513 6273 25547 6307
rect 25697 6273 25731 6307
rect 2973 6205 3007 6239
rect 7941 6205 7975 6239
rect 8309 6205 8343 6239
rect 11345 6205 11379 6239
rect 12357 6205 12391 6239
rect 19073 6205 19107 6239
rect 23673 6205 23707 6239
rect 6469 6137 6503 6171
rect 2513 6069 2547 6103
rect 5365 6069 5399 6103
rect 5549 6069 5583 6103
rect 5641 6069 5675 6103
rect 7665 6069 7699 6103
rect 9505 6069 9539 6103
rect 9689 6069 9723 6103
rect 10701 6069 10735 6103
rect 14657 6069 14691 6103
rect 20453 6069 20487 6103
rect 21557 6069 21591 6103
rect 25053 6069 25087 6103
rect 25145 6069 25179 6103
rect 4813 5865 4847 5899
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 14105 5865 14139 5899
rect 14933 5865 14967 5899
rect 23857 5865 23891 5899
rect 25789 5865 25823 5899
rect 6653 5797 6687 5831
rect 8217 5797 8251 5831
rect 16957 5797 16991 5831
rect 17693 5797 17727 5831
rect 25421 5797 25455 5831
rect 8125 5729 8159 5763
rect 15577 5729 15611 5763
rect 3065 5661 3099 5695
rect 5273 5661 5307 5695
rect 7858 5661 7892 5695
rect 10333 5661 10367 5695
rect 10517 5661 10551 5695
rect 10784 5661 10818 5695
rect 13921 5661 13955 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 15117 5661 15151 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 15485 5661 15519 5695
rect 17693 5661 17727 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 18429 5661 18463 5695
rect 20269 5661 20303 5695
rect 20545 5661 20579 5695
rect 20729 5661 20763 5695
rect 23765 5661 23799 5695
rect 24593 5661 24627 5695
rect 24685 5661 24719 5695
rect 24961 5661 24995 5695
rect 25053 5661 25087 5695
rect 25605 5661 25639 5695
rect 2881 5593 2915 5627
rect 4997 5593 5031 5627
rect 5181 5593 5215 5627
rect 5540 5593 5574 5627
rect 8585 5593 8619 5627
rect 10066 5593 10100 5627
rect 13737 5593 13771 5627
rect 15844 5593 15878 5627
rect 17233 5593 17267 5627
rect 17417 5593 17451 5627
rect 18061 5593 18095 5627
rect 20637 5593 20671 5627
rect 20996 5593 21030 5627
rect 23581 5593 23615 5627
rect 24041 5593 24075 5627
rect 24225 5593 24259 5627
rect 24777 5593 24811 5627
rect 25237 5593 25271 5627
rect 3249 5525 3283 5559
rect 6745 5525 6779 5559
rect 8769 5525 8803 5559
rect 11897 5525 11931 5559
rect 13553 5525 13587 5559
rect 17049 5525 17083 5559
rect 22109 5525 22143 5559
rect 23397 5525 23431 5559
rect 24409 5525 24443 5559
rect 4419 5321 4453 5355
rect 5549 5321 5583 5355
rect 5733 5321 5767 5355
rect 6577 5321 6611 5355
rect 6745 5321 6779 5355
rect 7849 5321 7883 5355
rect 15761 5321 15795 5355
rect 19533 5321 19567 5355
rect 24041 5321 24075 5355
rect 25513 5321 25547 5355
rect 25789 5321 25823 5355
rect 4629 5253 4663 5287
rect 6377 5253 6411 5287
rect 7481 5253 7515 5287
rect 7665 5253 7699 5287
rect 14013 5253 14047 5287
rect 14381 5253 14415 5287
rect 15025 5253 15059 5287
rect 20361 5253 20395 5287
rect 24378 5253 24412 5287
rect 1961 5185 1995 5219
rect 2145 5185 2179 5219
rect 2697 5185 2731 5219
rect 3913 5185 3947 5219
rect 4169 5185 4203 5219
rect 6101 5185 6135 5219
rect 9054 5185 9088 5219
rect 9321 5185 9355 5219
rect 13553 5185 13587 5219
rect 13645 5185 13679 5219
rect 13737 5185 13771 5219
rect 13921 5185 13955 5219
rect 14197 5185 14231 5219
rect 15209 5185 15243 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 16037 5185 16071 5219
rect 16129 5185 16163 5219
rect 16221 5185 16255 5219
rect 16405 5185 16439 5219
rect 18409 5185 18443 5219
rect 20177 5185 20211 5219
rect 20269 5185 20303 5219
rect 20545 5185 20579 5219
rect 21281 5185 21315 5219
rect 21373 5185 21407 5219
rect 21465 5185 21499 5219
rect 21649 5185 21683 5219
rect 21833 5185 21867 5219
rect 22089 5185 22123 5219
rect 23397 5185 23431 5219
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 23765 5185 23799 5219
rect 24133 5185 24167 5219
rect 25605 5185 25639 5219
rect 18153 5117 18187 5151
rect 21005 5117 21039 5151
rect 2053 5049 2087 5083
rect 2421 5049 2455 5083
rect 2789 5049 2823 5083
rect 4261 5049 4295 5083
rect 7941 5049 7975 5083
rect 2237 4981 2271 5015
rect 4445 4981 4479 5015
rect 5733 4981 5767 5015
rect 6561 4981 6595 5015
rect 13277 4981 13311 5015
rect 19993 4981 20027 5015
rect 23213 4981 23247 5015
rect 3525 4777 3559 4811
rect 8309 4777 8343 4811
rect 15117 4777 15151 4811
rect 15853 4777 15887 4811
rect 18061 4777 18095 4811
rect 18889 4777 18923 4811
rect 21649 4777 21683 4811
rect 21925 4777 21959 4811
rect 25789 4777 25823 4811
rect 2145 4641 2179 4675
rect 24409 4641 24443 4675
rect 2401 4573 2435 4607
rect 8217 4573 8251 4607
rect 8401 4573 8435 4607
rect 12541 4573 12575 4607
rect 12808 4573 12842 4607
rect 14381 4573 14415 4607
rect 14473 4573 14507 4607
rect 14565 4573 14599 4607
rect 14749 4573 14783 4607
rect 14933 4573 14967 4607
rect 16037 4573 16071 4607
rect 16405 4573 16439 4607
rect 18317 4573 18351 4607
rect 18429 4573 18463 4607
rect 18521 4573 18555 4607
rect 18705 4573 18739 4607
rect 19073 4573 19107 4607
rect 19441 4573 19475 4607
rect 21465 4573 21499 4607
rect 21741 4573 21775 4607
rect 23581 4573 23615 4607
rect 23765 4573 23799 4607
rect 23857 4573 23891 4607
rect 23949 4573 23983 4607
rect 16129 4505 16163 4539
rect 16221 4505 16255 4539
rect 19257 4505 19291 4539
rect 19625 4505 19659 4539
rect 21281 4505 21315 4539
rect 24225 4505 24259 4539
rect 24654 4505 24688 4539
rect 13921 4437 13955 4471
rect 14105 4437 14139 4471
rect 19625 4233 19659 4267
rect 16681 4165 16715 4199
rect 17049 4165 17083 4199
rect 20545 4165 20579 4199
rect 21281 4165 21315 4199
rect 21465 4165 21499 4199
rect 12900 4097 12934 4131
rect 14657 4097 14691 4131
rect 14749 4097 14783 4131
rect 14841 4097 14875 4131
rect 15025 4097 15059 4131
rect 15393 4097 15427 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 16037 4097 16071 4131
rect 16129 4097 16163 4131
rect 16221 4097 16255 4131
rect 16405 4097 16439 4131
rect 16865 4097 16899 4131
rect 17141 4097 17175 4131
rect 17325 4097 17359 4131
rect 17417 4097 17451 4131
rect 17509 4097 17543 4131
rect 18153 4097 18187 4131
rect 18420 4097 18454 4131
rect 19901 4097 19935 4131
rect 19993 4097 20027 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 20361 4097 20395 4131
rect 20637 4097 20671 4131
rect 20729 4097 20763 4131
rect 21833 4097 21867 4131
rect 22017 4097 22051 4131
rect 22109 4097 22143 4131
rect 22201 4097 22235 4131
rect 22937 4097 22971 4131
rect 23029 4097 23063 4131
rect 23121 4097 23155 4131
rect 23305 4097 23339 4131
rect 24613 4097 24647 4131
rect 24869 4097 24903 4131
rect 25237 4097 25271 4131
rect 25605 4097 25639 4131
rect 12633 4029 12667 4063
rect 21649 4029 21683 4063
rect 15853 3961 15887 3995
rect 19533 3961 19567 3995
rect 25421 3961 25455 3995
rect 25789 3961 25823 3995
rect 14013 3893 14047 3927
rect 14381 3893 14415 3927
rect 15117 3893 15151 3927
rect 17785 3893 17819 3927
rect 20913 3893 20947 3927
rect 22477 3893 22511 3927
rect 22661 3893 22695 3927
rect 23489 3893 23523 3927
rect 15485 3689 15519 3723
rect 18981 3689 19015 3723
rect 19257 3689 19291 3723
rect 23673 3689 23707 3723
rect 25053 3689 25087 3723
rect 18705 3621 18739 3655
rect 22109 3553 22143 3587
rect 22201 3553 22235 3587
rect 14105 3485 14139 3519
rect 15853 3485 15887 3519
rect 17325 3485 17359 3519
rect 19533 3485 19567 3519
rect 19625 3485 19659 3519
rect 19717 3485 19751 3519
rect 19901 3485 19935 3519
rect 19993 3485 20027 3519
rect 20177 3485 20211 3519
rect 20269 3485 20303 3519
rect 20385 3485 20419 3519
rect 22468 3485 22502 3519
rect 24041 3485 24075 3519
rect 24409 3485 24443 3519
rect 24593 3485 24627 3519
rect 24685 3485 24719 3519
rect 24777 3485 24811 3519
rect 25605 3485 25639 3519
rect 14372 3417 14406 3451
rect 16120 3417 16154 3451
rect 17592 3417 17626 3451
rect 18889 3417 18923 3451
rect 21842 3417 21876 3451
rect 23857 3417 23891 3451
rect 17233 3349 17267 3383
rect 20545 3349 20579 3383
rect 20729 3349 20763 3383
rect 23581 3349 23615 3383
rect 25789 3349 25823 3383
rect 15209 3145 15243 3179
rect 16681 3145 16715 3179
rect 17509 3145 17543 3179
rect 19809 3145 19843 3179
rect 20269 3145 20303 3179
rect 21465 3145 21499 3179
rect 21833 3145 21867 3179
rect 24041 3145 24075 3179
rect 24501 3145 24535 3179
rect 14004 3077 14038 3111
rect 15669 3077 15703 3111
rect 15853 3077 15887 3111
rect 17693 3077 17727 3111
rect 19104 3077 19138 3111
rect 20637 3077 20671 3111
rect 22928 3077 22962 3111
rect 24133 3077 24167 3111
rect 13737 3009 13771 3043
rect 15404 3009 15438 3043
rect 15577 3009 15611 3043
rect 16037 3009 16071 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 17141 3009 17175 3043
rect 17325 3009 17359 3043
rect 17877 3009 17911 3043
rect 19441 3009 19475 3043
rect 19625 3009 19659 3043
rect 20429 3009 20463 3043
rect 20545 3009 20579 3043
rect 20821 3009 20855 3043
rect 20913 3009 20947 3043
rect 21097 3009 21131 3043
rect 21189 3009 21223 3043
rect 21281 3009 21315 3043
rect 22109 3009 22143 3043
rect 22201 3009 22235 3043
rect 22293 3009 22327 3043
rect 22477 3009 22511 3043
rect 22661 3009 22695 3043
rect 24317 3009 24351 3043
rect 25605 3009 25639 3043
rect 19349 2941 19383 2975
rect 15117 2873 15151 2907
rect 17969 2805 18003 2839
rect 25789 2805 25823 2839
rect 10609 2601 10643 2635
rect 22017 2601 22051 2635
rect 19349 2533 19383 2567
rect 21557 2533 21591 2567
rect 22385 2533 22419 2567
rect 12633 2465 12667 2499
rect 10425 2397 10459 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 13553 2397 13587 2431
rect 13921 2397 13955 2431
rect 14565 2397 14599 2431
rect 15209 2397 15243 2431
rect 15853 2397 15887 2431
rect 16497 2397 16531 2431
rect 17141 2397 17175 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 18429 2397 18463 2431
rect 18613 2397 18647 2431
rect 19533 2397 19567 2431
rect 19901 2397 19935 2431
rect 20361 2397 20395 2431
rect 20729 2397 20763 2431
rect 21189 2397 21223 2431
rect 21833 2397 21867 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23305 2397 23339 2431
rect 23949 2397 23983 2431
rect 24869 2397 24903 2431
rect 18797 2329 18831 2363
rect 21373 2329 21407 2363
rect 11805 2261 11839 2295
rect 13369 2261 13403 2295
rect 13737 2261 13771 2295
rect 14381 2261 14415 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 16313 2261 16347 2295
rect 16957 2261 16991 2295
rect 17601 2261 17635 2295
rect 18153 2261 18187 2295
rect 19717 2261 19751 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
rect 22753 2261 22787 2295
rect 23489 2261 23523 2295
rect 24133 2261 24167 2295
rect 24685 2261 24719 2295
<< metal1 >>
rect 1104 27226 26220 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 26220 27226
rect 1104 27152 26220 27174
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 13081 27115 13139 27121
rect 13081 27112 13093 27115
rect 12952 27084 13093 27112
rect 12952 27072 12958 27084
rect 13081 27081 13093 27084
rect 13127 27081 13139 27115
rect 13081 27075 13139 27081
rect 13170 26936 13176 26988
rect 13228 26976 13234 26988
rect 13265 26979 13323 26985
rect 13265 26976 13277 26979
rect 13228 26948 13277 26976
rect 13228 26936 13234 26948
rect 13265 26945 13277 26948
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 1104 26682 26220 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 26220 26682
rect 1104 26608 26220 26630
rect 1104 26138 26220 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 26220 26138
rect 1104 26064 26220 26086
rect 1104 25594 26220 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 26220 25594
rect 1104 25520 26220 25542
rect 1104 25050 26220 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 26220 25050
rect 1104 24976 26220 24998
rect 9398 24760 9404 24812
rect 9456 24800 9462 24812
rect 11241 24803 11299 24809
rect 11241 24800 11253 24803
rect 9456 24772 11253 24800
rect 9456 24760 9462 24772
rect 11241 24769 11253 24772
rect 11287 24769 11299 24803
rect 11241 24763 11299 24769
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24800 11759 24803
rect 11882 24800 11888 24812
rect 11747 24772 11888 24800
rect 11747 24769 11759 24772
rect 11701 24763 11759 24769
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 12066 24809 12072 24812
rect 12060 24763 12072 24809
rect 12066 24760 12072 24763
rect 12124 24760 12130 24812
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 13964 24772 14381 24800
rect 13964 24760 13970 24772
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 21361 24803 21419 24809
rect 21361 24769 21373 24803
rect 21407 24800 21419 24803
rect 21726 24800 21732 24812
rect 21407 24772 21732 24800
rect 21407 24769 21419 24772
rect 21361 24763 21419 24769
rect 21726 24760 21732 24772
rect 21784 24760 21790 24812
rect 11790 24692 11796 24744
rect 11848 24692 11854 24744
rect 13354 24692 13360 24744
rect 13412 24732 13418 24744
rect 13817 24735 13875 24741
rect 13817 24732 13829 24735
rect 13412 24704 13829 24732
rect 13412 24692 13418 24704
rect 13817 24701 13829 24704
rect 13863 24701 13875 24735
rect 13817 24695 13875 24701
rect 10870 24624 10876 24676
rect 10928 24664 10934 24676
rect 11609 24667 11667 24673
rect 11609 24664 11621 24667
rect 10928 24636 11621 24664
rect 10928 24624 10934 24636
rect 11609 24633 11621 24636
rect 11655 24633 11667 24667
rect 11609 24627 11667 24633
rect 13170 24624 13176 24676
rect 13228 24624 13234 24676
rect 11054 24556 11060 24608
rect 11112 24556 11118 24608
rect 13262 24556 13268 24608
rect 13320 24556 13326 24608
rect 14274 24556 14280 24608
rect 14332 24556 14338 24608
rect 21174 24556 21180 24608
rect 21232 24556 21238 24608
rect 1104 24506 26220 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 26220 24506
rect 1104 24432 26220 24454
rect 13262 24392 13268 24404
rect 12084 24364 13268 24392
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11422 24188 11428 24200
rect 11379 24160 11428 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 11624 24120 11652 24151
rect 11698 24148 11704 24200
rect 11756 24188 11762 24200
rect 12084 24197 12112 24364
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 18417 24395 18475 24401
rect 18417 24392 18429 24395
rect 18156 24364 18429 24392
rect 12526 24324 12532 24336
rect 12176 24296 12532 24324
rect 12176 24265 12204 24296
rect 12526 24284 12532 24296
rect 12584 24284 12590 24336
rect 12161 24259 12219 24265
rect 12161 24225 12173 24259
rect 12207 24225 12219 24259
rect 18156 24256 18184 24364
rect 18417 24361 18429 24364
rect 18463 24361 18475 24395
rect 18417 24355 18475 24361
rect 12161 24219 12219 24225
rect 12268 24228 12673 24256
rect 11793 24191 11851 24197
rect 11793 24188 11805 24191
rect 11756 24160 11805 24188
rect 11756 24148 11762 24160
rect 11793 24157 11805 24160
rect 11839 24157 11851 24191
rect 11793 24151 11851 24157
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 11882 24120 11888 24132
rect 11624 24092 11888 24120
rect 11882 24080 11888 24092
rect 11940 24080 11946 24132
rect 12268 24064 12296 24228
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12400 24160 12541 24188
rect 12400 24148 12406 24160
rect 12529 24157 12541 24160
rect 12575 24157 12587 24191
rect 12645 24188 12673 24228
rect 18064 24228 18184 24256
rect 18417 24259 18475 24265
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 12645 24160 14105 24188
rect 12529 24151 12587 24157
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 16301 24191 16359 24197
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 17586 24188 17592 24200
rect 16531 24160 17592 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 12774 24123 12832 24129
rect 12774 24120 12786 24123
rect 12452 24092 12786 24120
rect 10689 24055 10747 24061
rect 10689 24021 10701 24055
rect 10735 24052 10747 24055
rect 10962 24052 10968 24064
rect 10735 24024 10968 24052
rect 10735 24021 10747 24024
rect 10689 24015 10747 24021
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12250 24052 12256 24064
rect 11747 24024 12256 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 12452 24061 12480 24092
rect 12774 24089 12786 24092
rect 12820 24089 12832 24123
rect 12774 24083 12832 24089
rect 13170 24080 13176 24132
rect 13228 24120 13234 24132
rect 14277 24123 14335 24129
rect 14277 24120 14289 24123
rect 13228 24092 14289 24120
rect 13228 24080 13234 24092
rect 14277 24089 14289 24092
rect 14323 24089 14335 24123
rect 16316 24120 16344 24151
rect 17586 24148 17592 24160
rect 17644 24148 17650 24200
rect 17885 24191 17943 24197
rect 17885 24157 17897 24191
rect 17931 24188 17943 24191
rect 18064 24188 18092 24228
rect 18417 24225 18429 24259
rect 18463 24225 18475 24259
rect 18417 24219 18475 24225
rect 18509 24259 18567 24265
rect 18509 24225 18521 24259
rect 18555 24256 18567 24259
rect 18969 24259 19027 24265
rect 18555 24228 18828 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 17931 24160 18092 24188
rect 17931 24157 17943 24160
rect 17885 24151 17943 24157
rect 18138 24148 18144 24200
rect 18196 24148 18202 24200
rect 18233 24123 18291 24129
rect 18233 24120 18245 24123
rect 16316 24092 18245 24120
rect 14277 24083 14335 24089
rect 18233 24089 18245 24092
rect 18279 24120 18291 24123
rect 18322 24120 18328 24132
rect 18279 24092 18328 24120
rect 18279 24089 18291 24092
rect 18233 24083 18291 24089
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 12437 24055 12495 24061
rect 12437 24021 12449 24055
rect 12483 24021 12495 24055
rect 12437 24015 12495 24021
rect 13354 24012 13360 24064
rect 13412 24052 13418 24064
rect 13909 24055 13967 24061
rect 13909 24052 13921 24055
rect 13412 24024 13921 24052
rect 13412 24012 13418 24024
rect 13909 24021 13921 24024
rect 13955 24021 13967 24055
rect 13909 24015 13967 24021
rect 14458 24012 14464 24064
rect 14516 24012 14522 24064
rect 16393 24055 16451 24061
rect 16393 24021 16405 24055
rect 16439 24052 16451 24055
rect 16574 24052 16580 24064
rect 16439 24024 16580 24052
rect 16439 24021 16451 24024
rect 16393 24015 16451 24021
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 16758 24012 16764 24064
rect 16816 24012 16822 24064
rect 17862 24012 17868 24064
rect 17920 24052 17926 24064
rect 18432 24052 18460 24219
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24157 18659 24191
rect 18601 24151 18659 24157
rect 17920 24024 18460 24052
rect 18616 24052 18644 24151
rect 18690 24148 18696 24200
rect 18748 24148 18754 24200
rect 18800 24197 18828 24228
rect 18969 24225 18981 24259
rect 19015 24256 19027 24259
rect 19242 24256 19248 24268
rect 19015 24228 19248 24256
rect 19015 24225 19027 24228
rect 18969 24219 19027 24225
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 18785 24191 18843 24197
rect 18785 24157 18797 24191
rect 18831 24188 18843 24191
rect 19702 24188 19708 24200
rect 18831 24160 19708 24188
rect 18831 24157 18843 24160
rect 18785 24151 18843 24157
rect 19702 24148 19708 24160
rect 19760 24148 19766 24200
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24188 21603 24191
rect 23017 24191 23075 24197
rect 23017 24188 23029 24191
rect 21591 24160 23029 24188
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 23017 24157 23029 24160
rect 23063 24188 23075 24191
rect 23382 24188 23388 24200
rect 23063 24160 23388 24188
rect 23063 24157 23075 24160
rect 23017 24151 23075 24157
rect 23382 24148 23388 24160
rect 23440 24148 23446 24200
rect 19610 24120 19616 24132
rect 18892 24092 19616 24120
rect 18892 24052 18920 24092
rect 19610 24080 19616 24092
rect 19668 24080 19674 24132
rect 21082 24080 21088 24132
rect 21140 24120 21146 24132
rect 21278 24123 21336 24129
rect 21278 24120 21290 24123
rect 21140 24092 21290 24120
rect 21140 24080 21146 24092
rect 21278 24089 21290 24092
rect 21324 24089 21336 24123
rect 21278 24083 21336 24089
rect 21450 24080 21456 24132
rect 21508 24120 21514 24132
rect 22750 24123 22808 24129
rect 22750 24120 22762 24123
rect 21508 24092 22762 24120
rect 21508 24080 21514 24092
rect 22750 24089 22762 24092
rect 22796 24089 22808 24123
rect 22750 24083 22808 24089
rect 18616 24024 18920 24052
rect 18969 24055 19027 24061
rect 17920 24012 17926 24024
rect 18969 24021 18981 24055
rect 19015 24052 19027 24055
rect 19426 24052 19432 24064
rect 19015 24024 19432 24052
rect 19015 24021 19027 24024
rect 18969 24015 19027 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 20162 24012 20168 24064
rect 20220 24012 20226 24064
rect 21637 24055 21695 24061
rect 21637 24021 21649 24055
rect 21683 24052 21695 24055
rect 21726 24052 21732 24064
rect 21683 24024 21732 24052
rect 21683 24021 21695 24024
rect 21637 24015 21695 24021
rect 21726 24012 21732 24024
rect 21784 24012 21790 24064
rect 1104 23962 26220 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 26220 23962
rect 1104 23888 26220 23910
rect 9398 23848 9404 23860
rect 8772 23820 9404 23848
rect 8772 23789 8800 23820
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 11790 23808 11796 23860
rect 11848 23808 11854 23860
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 12434 23848 12440 23860
rect 11940 23820 12440 23848
rect 11940 23808 11946 23820
rect 12434 23808 12440 23820
rect 12492 23848 12498 23860
rect 12897 23851 12955 23857
rect 12897 23848 12909 23851
rect 12492 23820 12909 23848
rect 12492 23808 12498 23820
rect 12897 23817 12909 23820
rect 12943 23817 12955 23851
rect 12897 23811 12955 23817
rect 21361 23851 21419 23857
rect 21361 23817 21373 23851
rect 21407 23848 21419 23851
rect 21450 23848 21456 23860
rect 21407 23820 21456 23848
rect 21407 23817 21419 23820
rect 21361 23811 21419 23817
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 8757 23783 8815 23789
rect 8757 23749 8769 23783
rect 8803 23749 8815 23783
rect 11808 23780 11836 23808
rect 12342 23780 12348 23792
rect 8757 23743 8815 23749
rect 10796 23752 12348 23780
rect 10502 23672 10508 23724
rect 10560 23721 10566 23724
rect 10796 23721 10824 23752
rect 10560 23675 10572 23721
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23681 10839 23715
rect 10781 23675 10839 23681
rect 10560 23672 10566 23675
rect 10870 23672 10876 23724
rect 10928 23672 10934 23724
rect 10962 23672 10968 23724
rect 11020 23672 11026 23724
rect 11532 23721 11560 23752
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 13633 23783 13691 23789
rect 13633 23749 13645 23783
rect 13679 23780 13691 23783
rect 14458 23780 14464 23792
rect 13679 23752 14464 23780
rect 13679 23749 13691 23752
rect 13633 23743 13691 23749
rect 14458 23740 14464 23752
rect 14516 23740 14522 23792
rect 16482 23740 16488 23792
rect 16540 23780 16546 23792
rect 18138 23780 18144 23792
rect 16540 23752 18144 23780
rect 16540 23740 16546 23752
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11784 23715 11842 23721
rect 11784 23681 11796 23715
rect 11830 23712 11842 23715
rect 12158 23712 12164 23724
rect 11830 23684 12164 23712
rect 11830 23681 11842 23684
rect 11784 23675 11842 23681
rect 12158 23672 12164 23684
rect 12216 23672 12222 23724
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 13265 23715 13323 23721
rect 13265 23712 13277 23715
rect 12584 23684 13277 23712
rect 12584 23672 12590 23684
rect 13265 23681 13277 23684
rect 13311 23712 13323 23715
rect 13998 23712 14004 23724
rect 13311 23684 14004 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 14550 23672 14556 23724
rect 14608 23672 14614 23724
rect 14734 23672 14740 23724
rect 14792 23672 14798 23724
rect 17793 23715 17851 23721
rect 17793 23681 17805 23715
rect 17839 23712 17851 23715
rect 17954 23712 17960 23724
rect 17839 23684 17960 23712
rect 17839 23681 17851 23684
rect 17793 23675 17851 23681
rect 17954 23672 17960 23684
rect 18012 23672 18018 23724
rect 18064 23721 18092 23752
rect 18138 23740 18144 23752
rect 18196 23740 18202 23792
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23712 18107 23715
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 18095 23684 19073 23712
rect 18095 23681 18107 23684
rect 18049 23675 18107 23681
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19150 23672 19156 23724
rect 19208 23712 19214 23724
rect 19317 23715 19375 23721
rect 19317 23712 19329 23715
rect 19208 23684 19329 23712
rect 19208 23672 19214 23684
rect 19317 23681 19329 23684
rect 19363 23681 19375 23715
rect 19317 23675 19375 23681
rect 20622 23672 20628 23724
rect 20680 23712 20686 23724
rect 20901 23715 20959 23721
rect 20901 23712 20913 23715
rect 20680 23684 20913 23712
rect 20680 23672 20686 23684
rect 20901 23681 20913 23684
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23613 4951 23647
rect 4893 23607 4951 23613
rect 4614 23536 4620 23588
rect 4672 23576 4678 23588
rect 4908 23576 4936 23607
rect 5166 23604 5172 23656
rect 5224 23604 5230 23656
rect 5258 23604 5264 23656
rect 5316 23604 5322 23656
rect 5378 23647 5436 23653
rect 5378 23613 5390 23647
rect 5424 23644 5436 23647
rect 5994 23644 6000 23656
rect 5424 23616 6000 23644
rect 5424 23613 5436 23616
rect 5378 23607 5436 23613
rect 5994 23604 6000 23616
rect 6052 23604 6058 23656
rect 11146 23604 11152 23656
rect 11204 23604 11210 23656
rect 11238 23604 11244 23656
rect 11296 23604 11302 23656
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23644 13231 23647
rect 13354 23644 13360 23656
rect 13219 23616 13360 23644
rect 13219 23613 13231 23616
rect 13173 23607 13231 23613
rect 13354 23604 13360 23616
rect 13412 23604 13418 23656
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14277 23607 14335 23613
rect 13372 23576 13400 23604
rect 14292 23576 14320 23607
rect 16206 23604 16212 23656
rect 16264 23604 16270 23656
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23613 18199 23647
rect 18141 23607 18199 23613
rect 20809 23647 20867 23653
rect 20809 23613 20821 23647
rect 20855 23644 20867 23647
rect 21174 23644 21180 23656
rect 20855 23616 21180 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 4672 23548 5488 23576
rect 13372 23548 14320 23576
rect 4672 23536 4678 23548
rect 5460 23520 5488 23548
rect 5442 23468 5448 23520
rect 5500 23468 5506 23520
rect 5534 23468 5540 23520
rect 5592 23468 5598 23520
rect 8662 23468 8668 23520
rect 8720 23468 8726 23520
rect 11330 23468 11336 23520
rect 11388 23468 11394 23520
rect 12986 23468 12992 23520
rect 13044 23468 13050 23520
rect 13078 23468 13084 23520
rect 13136 23508 13142 23520
rect 13725 23511 13783 23517
rect 13725 23508 13737 23511
rect 13136 23480 13737 23508
rect 13136 23468 13142 23480
rect 13725 23477 13737 23480
rect 13771 23477 13783 23511
rect 13725 23471 13783 23477
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14737 23511 14795 23517
rect 14737 23508 14749 23511
rect 13872 23480 14749 23508
rect 13872 23468 13878 23480
rect 14737 23477 14749 23480
rect 14783 23477 14795 23511
rect 14737 23471 14795 23477
rect 15562 23468 15568 23520
rect 15620 23508 15626 23520
rect 15657 23511 15715 23517
rect 15657 23508 15669 23511
rect 15620 23480 15669 23508
rect 15620 23468 15626 23480
rect 15657 23477 15669 23480
rect 15703 23477 15715 23511
rect 15657 23471 15715 23477
rect 16666 23468 16672 23520
rect 16724 23508 16730 23520
rect 17770 23508 17776 23520
rect 16724 23480 17776 23508
rect 16724 23468 16730 23480
rect 17770 23468 17776 23480
rect 17828 23508 17834 23520
rect 18156 23508 18184 23607
rect 21174 23604 21180 23616
rect 21232 23604 21238 23656
rect 17828 23480 18184 23508
rect 17828 23468 17834 23480
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 18785 23511 18843 23517
rect 18785 23508 18797 23511
rect 18748 23480 18797 23508
rect 18748 23468 18754 23480
rect 18785 23477 18797 23480
rect 18831 23477 18843 23511
rect 18785 23471 18843 23477
rect 20254 23468 20260 23520
rect 20312 23508 20318 23520
rect 20441 23511 20499 23517
rect 20441 23508 20453 23511
rect 20312 23480 20453 23508
rect 20312 23468 20318 23480
rect 20441 23477 20453 23480
rect 20487 23477 20499 23511
rect 20441 23471 20499 23477
rect 1104 23418 26220 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 26220 23418
rect 1104 23344 26220 23366
rect 5258 23304 5264 23316
rect 5006 23276 5264 23304
rect 3602 23196 3608 23248
rect 3660 23196 3666 23248
rect 3694 23196 3700 23248
rect 3752 23236 3758 23248
rect 5006 23236 5034 23276
rect 5258 23264 5264 23276
rect 5316 23304 5322 23316
rect 8478 23304 8484 23316
rect 5316 23276 8484 23304
rect 5316 23264 5322 23276
rect 8478 23264 8484 23276
rect 8536 23264 8542 23316
rect 10502 23264 10508 23316
rect 10560 23264 10566 23316
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 11072 23276 11345 23304
rect 3752 23208 5034 23236
rect 3752 23196 3758 23208
rect 3234 23128 3240 23180
rect 3292 23168 3298 23180
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 3292 23140 4261 23168
rect 3292 23128 3298 23140
rect 4249 23137 4261 23140
rect 4295 23168 4307 23171
rect 4430 23168 4436 23180
rect 4295 23140 4436 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 4632 23177 4660 23208
rect 4617 23171 4675 23177
rect 4617 23137 4629 23171
rect 4663 23137 4675 23171
rect 4617 23131 4675 23137
rect 4706 23128 4712 23180
rect 4764 23177 4770 23180
rect 4764 23171 4792 23177
rect 4780 23137 4792 23171
rect 4764 23131 4792 23137
rect 10689 23171 10747 23177
rect 10689 23137 10701 23171
rect 10735 23168 10747 23171
rect 10870 23168 10876 23180
rect 10735 23140 10876 23168
rect 10735 23137 10747 23140
rect 10689 23131 10747 23137
rect 4764 23128 4770 23131
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 1946 23060 1952 23112
rect 2004 23100 2010 23112
rect 2225 23103 2283 23109
rect 2225 23100 2237 23103
rect 2004 23072 2237 23100
rect 2004 23060 2010 23072
rect 2225 23069 2237 23072
rect 2271 23069 2283 23103
rect 4985 23103 5043 23109
rect 4985 23100 4997 23103
rect 2225 23063 2283 23069
rect 4632 23072 4997 23100
rect 4632 23044 4660 23072
rect 4985 23069 4997 23072
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 5252 23103 5310 23109
rect 5252 23069 5264 23103
rect 5298 23100 5310 23103
rect 5534 23100 5540 23112
rect 5298 23072 5540 23100
rect 5298 23069 5310 23072
rect 5252 23063 5310 23069
rect 5534 23060 5540 23072
rect 5592 23060 5598 23112
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23100 7251 23103
rect 8294 23100 8300 23112
rect 7239 23072 8300 23100
rect 7239 23069 7251 23072
rect 7193 23063 7251 23069
rect 8294 23060 8300 23072
rect 8352 23100 8358 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8352 23072 8953 23100
rect 8352 23060 8358 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23100 10839 23103
rect 11072 23100 11100 23276
rect 11333 23273 11345 23276
rect 11379 23304 11391 23307
rect 11698 23304 11704 23316
rect 11379 23276 11704 23304
rect 11379 23273 11391 23276
rect 11333 23267 11391 23273
rect 11698 23264 11704 23276
rect 11756 23304 11762 23316
rect 11974 23304 11980 23316
rect 11756 23276 11980 23304
rect 11756 23264 11762 23276
rect 11974 23264 11980 23276
rect 12032 23264 12038 23316
rect 12158 23264 12164 23316
rect 12216 23264 12222 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 13265 23307 13323 23313
rect 13265 23304 13277 23307
rect 12492 23276 13277 23304
rect 12492 23264 12498 23276
rect 13265 23273 13277 23276
rect 13311 23304 13323 23307
rect 13722 23304 13728 23316
rect 13311 23276 13728 23304
rect 13311 23273 13323 23276
rect 13265 23267 13323 23273
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 13817 23307 13875 23313
rect 13817 23273 13829 23307
rect 13863 23304 13875 23307
rect 13998 23304 14004 23316
rect 13863 23276 14004 23304
rect 13863 23273 13875 23276
rect 13817 23267 13875 23273
rect 13998 23264 14004 23276
rect 14056 23264 14062 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 16816 23276 17816 23304
rect 16816 23264 16822 23276
rect 11422 23236 11428 23248
rect 11256 23208 11428 23236
rect 11256 23109 11284 23208
rect 11422 23196 11428 23208
rect 11480 23236 11486 23248
rect 11606 23236 11612 23248
rect 11480 23208 11612 23236
rect 11480 23196 11486 23208
rect 11606 23196 11612 23208
rect 11664 23196 11670 23248
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 12253 23239 12311 23245
rect 12253 23236 12265 23239
rect 12124 23208 12265 23236
rect 12124 23196 12130 23208
rect 12253 23205 12265 23208
rect 12299 23205 12311 23239
rect 12253 23199 12311 23205
rect 12529 23239 12587 23245
rect 12529 23205 12541 23239
rect 12575 23236 12587 23239
rect 14642 23236 14648 23248
rect 12575 23208 14648 23236
rect 12575 23205 12587 23208
rect 12529 23199 12587 23205
rect 14642 23196 14648 23208
rect 14700 23196 14706 23248
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 11388 23140 11529 23168
rect 11388 23128 11394 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 13078 23168 13084 23180
rect 11517 23131 11575 23137
rect 12452 23140 13084 23168
rect 10827 23072 11100 23100
rect 11241 23103 11299 23109
rect 10827 23069 10839 23072
rect 10781 23063 10839 23069
rect 11241 23069 11253 23103
rect 11287 23069 11299 23103
rect 11241 23063 11299 23069
rect 11433 23097 11491 23103
rect 11433 23063 11445 23097
rect 11479 23094 11491 23097
rect 11479 23066 11560 23094
rect 11479 23063 11491 23066
rect 2498 23041 2504 23044
rect 2492 22995 2504 23041
rect 2498 22992 2504 22995
rect 2556 22992 2562 23044
rect 4614 22992 4620 23044
rect 4672 22992 4678 23044
rect 5166 23032 5172 23044
rect 4816 23004 5172 23032
rect 2590 22924 2596 22976
rect 2648 22964 2654 22976
rect 4525 22967 4583 22973
rect 4525 22964 4537 22967
rect 2648 22936 4537 22964
rect 2648 22924 2654 22936
rect 4525 22933 4537 22936
rect 4571 22964 4583 22967
rect 4816 22964 4844 23004
rect 5166 22992 5172 23004
rect 5224 22992 5230 23044
rect 7006 22992 7012 23044
rect 7064 23032 7070 23044
rect 7438 23035 7496 23041
rect 7438 23032 7450 23035
rect 7064 23004 7450 23032
rect 7064 22992 7070 23004
rect 7438 23001 7450 23004
rect 7484 23001 7496 23035
rect 7438 22995 7496 23001
rect 8754 22992 8760 23044
rect 8812 23032 8818 23044
rect 9186 23035 9244 23041
rect 9186 23032 9198 23035
rect 8812 23004 9198 23032
rect 8812 22992 8818 23004
rect 9186 23001 9198 23004
rect 9232 23001 9244 23035
rect 9186 22995 9244 23001
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 11146 22992 11152 23044
rect 11204 22992 11210 23044
rect 4571 22936 4844 22964
rect 4571 22933 4583 22936
rect 4525 22927 4583 22933
rect 4890 22924 4896 22976
rect 4948 22924 4954 22976
rect 6362 22924 6368 22976
rect 6420 22924 6426 22976
rect 6638 22924 6644 22976
rect 6696 22964 6702 22976
rect 8573 22967 8631 22973
rect 8573 22964 8585 22967
rect 6696 22936 8585 22964
rect 6696 22924 6702 22936
rect 8573 22933 8585 22936
rect 8619 22964 8631 22967
rect 9030 22964 9036 22976
rect 8619 22936 9036 22964
rect 8619 22933 8631 22936
rect 8573 22927 8631 22933
rect 9030 22924 9036 22936
rect 9088 22924 9094 22976
rect 10321 22967 10379 22973
rect 10321 22933 10333 22967
rect 10367 22964 10379 22967
rect 11256 22964 11284 23063
rect 11433 23057 11491 23063
rect 10367 22936 11284 22964
rect 11532 22964 11560 23066
rect 12066 23060 12072 23112
rect 12124 23100 12130 23112
rect 12342 23100 12348 23112
rect 12124 23072 12348 23100
rect 12124 23060 12130 23072
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12452 23109 12480 23140
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 13814 23168 13820 23180
rect 13280 23140 13820 23168
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12526 23060 12532 23112
rect 12584 23100 12590 23112
rect 12621 23103 12679 23109
rect 12621 23100 12633 23103
rect 12584 23072 12633 23100
rect 12584 23060 12590 23072
rect 12621 23069 12633 23072
rect 12667 23069 12679 23103
rect 12621 23063 12679 23069
rect 12710 23060 12716 23112
rect 12768 23060 12774 23112
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 12986 23100 12992 23112
rect 12943 23072 12992 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 12986 23060 12992 23072
rect 13044 23060 13050 23112
rect 13280 23109 13308 23140
rect 13814 23128 13820 23140
rect 13872 23128 13878 23180
rect 16482 23168 16488 23180
rect 15672 23140 16488 23168
rect 15672 23112 15700 23140
rect 16482 23128 16488 23140
rect 16540 23128 16546 23180
rect 17788 23168 17816 23276
rect 18524 23276 18705 23304
rect 18524 23177 18552 23276
rect 18693 23273 18705 23276
rect 18739 23273 18751 23307
rect 18693 23267 18751 23273
rect 19150 23264 19156 23316
rect 19208 23304 19214 23316
rect 19245 23307 19303 23313
rect 19245 23304 19257 23307
rect 19208 23276 19257 23304
rect 19208 23264 19214 23276
rect 19245 23273 19257 23276
rect 19291 23273 19303 23307
rect 19245 23267 19303 23273
rect 19610 23264 19616 23316
rect 19668 23304 19674 23316
rect 19668 23276 20392 23304
rect 19668 23264 19674 23276
rect 19702 23196 19708 23248
rect 19760 23236 19766 23248
rect 19981 23239 20039 23245
rect 19981 23236 19993 23239
rect 19760 23208 19993 23236
rect 19760 23196 19766 23208
rect 19981 23205 19993 23208
rect 20027 23205 20039 23239
rect 20364 23236 20392 23276
rect 21082 23264 21088 23316
rect 21140 23264 21146 23316
rect 21542 23304 21548 23316
rect 21192 23276 21548 23304
rect 21192 23236 21220 23276
rect 21542 23264 21548 23276
rect 21600 23264 21606 23316
rect 20364 23208 21220 23236
rect 19981 23199 20039 23205
rect 21266 23196 21272 23248
rect 21324 23236 21330 23248
rect 21324 23208 22140 23236
rect 21324 23196 21330 23208
rect 18509 23171 18567 23177
rect 18509 23168 18521 23171
rect 17788 23140 18521 23168
rect 18509 23137 18521 23140
rect 18555 23137 18567 23171
rect 18785 23171 18843 23177
rect 18785 23168 18797 23171
rect 18509 23131 18567 23137
rect 18616 23140 18797 23168
rect 13265 23103 13323 23109
rect 13265 23069 13277 23103
rect 13311 23069 13323 23103
rect 13265 23063 13323 23069
rect 13354 23060 13360 23112
rect 13412 23060 13418 23112
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 13909 23103 13967 23109
rect 13909 23069 13921 23103
rect 13955 23069 13967 23103
rect 13909 23063 13967 23069
rect 15401 23103 15459 23109
rect 15401 23069 15413 23103
rect 15447 23100 15459 23103
rect 15562 23100 15568 23112
rect 15447 23072 15568 23100
rect 15447 23069 15459 23072
rect 15401 23063 15459 23069
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 13924 23032 13952 23063
rect 15562 23060 15568 23072
rect 15620 23060 15626 23112
rect 15654 23060 15660 23112
rect 15712 23060 15718 23112
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 13228 23004 13952 23032
rect 13228 22992 13234 23004
rect 13354 22964 13360 22976
rect 11532 22936 13360 22964
rect 10367 22933 10379 22936
rect 10321 22927 10379 22933
rect 13354 22924 13360 22936
rect 13412 22924 13418 22976
rect 13633 22967 13691 22973
rect 13633 22933 13645 22967
rect 13679 22964 13691 22967
rect 13722 22964 13728 22976
rect 13679 22936 13728 22964
rect 13679 22933 13691 22936
rect 13633 22927 13691 22933
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 14277 22967 14335 22973
rect 14277 22933 14289 22967
rect 14323 22964 14335 22967
rect 14550 22964 14556 22976
rect 14323 22936 14556 22964
rect 14323 22933 14335 22936
rect 14277 22927 14335 22933
rect 14550 22924 14556 22936
rect 14608 22964 14614 22976
rect 15764 22964 15792 23063
rect 16574 23060 16580 23112
rect 16632 23100 16638 23112
rect 16741 23103 16799 23109
rect 16741 23100 16753 23103
rect 16632 23072 16753 23100
rect 16632 23060 16638 23072
rect 16741 23069 16753 23072
rect 16787 23069 16799 23103
rect 16741 23063 16799 23069
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 18616 23100 18644 23140
rect 18785 23137 18797 23140
rect 18831 23168 18843 23171
rect 19150 23168 19156 23180
rect 18831 23140 19156 23168
rect 18831 23137 18843 23140
rect 18785 23131 18843 23137
rect 19150 23128 19156 23140
rect 19208 23128 19214 23180
rect 20530 23168 20536 23180
rect 19720 23140 20536 23168
rect 17828 23072 18644 23100
rect 18693 23103 18751 23109
rect 17828 23060 17834 23072
rect 18693 23069 18705 23103
rect 18739 23100 18751 23103
rect 18966 23100 18972 23112
rect 18739 23072 18972 23100
rect 18739 23069 18751 23072
rect 18693 23063 18751 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 19720 23109 19748 23140
rect 20530 23128 20536 23140
rect 20588 23128 20594 23180
rect 20990 23168 20996 23180
rect 20916 23140 20996 23168
rect 19521 23103 19579 23109
rect 19521 23069 19533 23103
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 19705 23103 19763 23109
rect 19705 23069 19717 23103
rect 19751 23069 19763 23103
rect 19705 23063 19763 23069
rect 18598 23032 18604 23044
rect 17880 23004 18604 23032
rect 14608 22936 15792 22964
rect 14608 22924 14614 22936
rect 16022 22924 16028 22976
rect 16080 22964 16086 22976
rect 16393 22967 16451 22973
rect 16393 22964 16405 22967
rect 16080 22936 16405 22964
rect 16080 22924 16086 22936
rect 16393 22933 16405 22936
rect 16439 22933 16451 22967
rect 16393 22927 16451 22933
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 17880 22973 17908 23004
rect 18598 22992 18604 23004
rect 18656 22992 18662 23044
rect 17865 22967 17923 22973
rect 17865 22964 17877 22967
rect 17092 22936 17877 22964
rect 17092 22924 17098 22936
rect 17865 22933 17877 22936
rect 17911 22933 17923 22967
rect 17865 22927 17923 22933
rect 17954 22924 17960 22976
rect 18012 22924 18018 22976
rect 19058 22924 19064 22976
rect 19116 22924 19122 22976
rect 19444 22964 19472 23060
rect 19536 23032 19564 23063
rect 19794 23060 19800 23112
rect 19852 23060 19858 23112
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23069 20039 23103
rect 19981 23063 20039 23069
rect 19996 23032 20024 23063
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 20916 23109 20944 23140
rect 20990 23128 20996 23140
rect 21048 23168 21054 23180
rect 21729 23171 21787 23177
rect 21729 23168 21741 23171
rect 21048 23140 21741 23168
rect 21048 23128 21054 23140
rect 21729 23137 21741 23140
rect 21775 23137 21787 23171
rect 21729 23131 21787 23137
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20220 23072 20453 23100
rect 20220 23060 20226 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20901 23103 20959 23109
rect 20901 23069 20913 23103
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 21174 23060 21180 23112
rect 21232 23060 21238 23112
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21545 23103 21603 23109
rect 21545 23100 21557 23103
rect 21324 23072 21557 23100
rect 21324 23060 21330 23072
rect 21545 23069 21557 23072
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21634 23060 21640 23112
rect 21692 23060 21698 23112
rect 21818 23060 21824 23112
rect 21876 23060 21882 23112
rect 22112 23109 22140 23208
rect 22186 23196 22192 23248
rect 22244 23236 22250 23248
rect 25685 23239 25743 23245
rect 25685 23236 25697 23239
rect 22244 23208 25697 23236
rect 22244 23196 22250 23208
rect 25685 23205 25697 23208
rect 25731 23205 25743 23239
rect 25685 23199 25743 23205
rect 21913 23103 21971 23109
rect 21913 23069 21925 23103
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 20254 23032 20260 23044
rect 19536 23004 20260 23032
rect 20254 22992 20260 23004
rect 20312 22992 20318 23044
rect 20622 23041 20628 23044
rect 20579 23035 20628 23041
rect 20579 23032 20591 23035
rect 20364 23004 20591 23032
rect 20364 22964 20392 23004
rect 20579 23001 20591 23004
rect 20625 23001 20628 23035
rect 20579 22995 20628 23001
rect 20622 22992 20628 22995
rect 20680 22992 20686 23044
rect 20717 23035 20775 23041
rect 20717 23001 20729 23035
rect 20763 23001 20775 23035
rect 20717 22995 20775 23001
rect 19444 22936 20392 22964
rect 20732 22964 20760 22995
rect 20806 22992 20812 23044
rect 20864 22992 20870 23044
rect 21192 23032 21220 23060
rect 21361 23035 21419 23041
rect 21361 23032 21373 23035
rect 21192 23004 21373 23032
rect 21361 23001 21373 23004
rect 21407 23001 21419 23035
rect 21361 22995 21419 23001
rect 21726 22992 21732 23044
rect 21784 23032 21790 23044
rect 21928 23032 21956 23063
rect 25222 23060 25228 23112
rect 25280 23060 25286 23112
rect 25866 23060 25872 23112
rect 25924 23060 25930 23112
rect 21784 23004 21956 23032
rect 21784 22992 21790 23004
rect 21174 22964 21180 22976
rect 20732 22936 21180 22964
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 21910 22924 21916 22976
rect 21968 22924 21974 22976
rect 25409 22967 25467 22973
rect 25409 22933 25421 22967
rect 25455 22964 25467 22967
rect 25590 22964 25596 22976
rect 25455 22936 25596 22964
rect 25455 22933 25467 22936
rect 25409 22927 25467 22933
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 1104 22874 26220 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 26220 22874
rect 1104 22800 26220 22822
rect 2498 22720 2504 22772
rect 2556 22720 2562 22772
rect 2590 22720 2596 22772
rect 2648 22760 2654 22772
rect 2869 22763 2927 22769
rect 2869 22760 2881 22763
rect 2648 22732 2881 22760
rect 2648 22720 2654 22732
rect 2869 22729 2881 22732
rect 2915 22729 2927 22763
rect 4982 22760 4988 22772
rect 2869 22723 2927 22729
rect 4172 22732 4988 22760
rect 4172 22701 4200 22732
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 5258 22720 5264 22772
rect 5316 22760 5322 22772
rect 5316 22732 6776 22760
rect 5316 22720 5322 22732
rect 4157 22695 4215 22701
rect 4157 22661 4169 22695
rect 4203 22661 4215 22695
rect 4357 22695 4415 22701
rect 4357 22692 4369 22695
rect 4157 22655 4215 22661
rect 4264 22664 4369 22692
rect 2660 22627 2718 22633
rect 2660 22593 2672 22627
rect 2706 22624 2718 22627
rect 2706 22596 3280 22624
rect 2706 22593 2718 22596
rect 2660 22587 2718 22593
rect 2774 22516 2780 22568
rect 2832 22516 2838 22568
rect 3142 22516 3148 22568
rect 3200 22516 3206 22568
rect 3252 22565 3280 22596
rect 3602 22584 3608 22636
rect 3660 22584 3666 22636
rect 4264 22624 4292 22664
rect 4357 22661 4369 22664
rect 4403 22661 4415 22695
rect 4357 22655 4415 22661
rect 4798 22652 4804 22704
rect 4856 22652 4862 22704
rect 6638 22692 6644 22704
rect 6564 22664 6644 22692
rect 3804 22596 4292 22624
rect 4816 22622 4844 22652
rect 6564 22633 6592 22664
rect 6638 22652 6644 22664
rect 6696 22652 6702 22704
rect 6748 22692 6776 22732
rect 7006 22720 7012 22772
rect 7064 22720 7070 22772
rect 7116 22732 8616 22760
rect 7116 22692 7144 22732
rect 6748 22664 7144 22692
rect 7285 22695 7343 22701
rect 7285 22661 7297 22695
rect 7331 22692 7343 22695
rect 7926 22692 7932 22704
rect 7331 22664 7932 22692
rect 7331 22661 7343 22664
rect 7285 22655 7343 22661
rect 7926 22652 7932 22664
rect 7984 22652 7990 22704
rect 8588 22636 8616 22732
rect 11606 22720 11612 22772
rect 11664 22760 11670 22772
rect 13170 22760 13176 22772
rect 11664 22732 13176 22760
rect 11664 22720 11670 22732
rect 13170 22720 13176 22732
rect 13228 22720 13234 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14792 22732 14933 22760
rect 14792 22720 14798 22732
rect 14921 22729 14933 22732
rect 14967 22729 14979 22763
rect 14921 22723 14979 22729
rect 15749 22763 15807 22769
rect 15749 22729 15761 22763
rect 15795 22760 15807 22763
rect 16206 22760 16212 22772
rect 15795 22732 16212 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 17865 22763 17923 22769
rect 17865 22760 17877 22763
rect 17144 22732 17877 22760
rect 8662 22652 8668 22704
rect 8720 22692 8726 22704
rect 8757 22695 8815 22701
rect 8757 22692 8769 22695
rect 8720 22664 8769 22692
rect 8720 22652 8726 22664
rect 8757 22661 8769 22664
rect 8803 22661 8815 22695
rect 8757 22655 8815 22661
rect 12161 22695 12219 22701
rect 12161 22661 12173 22695
rect 12207 22692 12219 22695
rect 12434 22692 12440 22704
rect 12207 22664 12440 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 12434 22652 12440 22664
rect 12492 22652 12498 22704
rect 13808 22695 13866 22701
rect 13808 22661 13820 22695
rect 13854 22692 13866 22695
rect 13906 22692 13912 22704
rect 13854 22664 13912 22692
rect 13854 22661 13866 22664
rect 13808 22655 13866 22661
rect 13906 22652 13912 22664
rect 13964 22652 13970 22704
rect 17144 22701 17172 22732
rect 17865 22729 17877 22732
rect 17911 22729 17923 22763
rect 17865 22723 17923 22729
rect 18046 22720 18052 22772
rect 18104 22760 18110 22772
rect 18141 22763 18199 22769
rect 18141 22760 18153 22763
rect 18104 22732 18153 22760
rect 18104 22720 18110 22732
rect 18141 22729 18153 22732
rect 18187 22729 18199 22763
rect 20651 22763 20709 22769
rect 18141 22723 18199 22729
rect 19536 22732 20208 22760
rect 17129 22695 17187 22701
rect 17129 22692 17141 22695
rect 16224 22664 17141 22692
rect 4884 22627 4942 22633
rect 4884 22622 4896 22627
rect 3804 22568 3832 22596
rect 4816 22594 4896 22622
rect 4884 22593 4896 22594
rect 4930 22593 4942 22627
rect 4884 22587 4942 22593
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7834 22624 7840 22636
rect 7423 22596 7840 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 8478 22584 8484 22636
rect 8536 22584 8542 22636
rect 8570 22584 8576 22636
rect 8628 22584 8634 22636
rect 11333 22627 11391 22633
rect 11333 22593 11345 22627
rect 11379 22593 11391 22627
rect 11333 22587 11391 22593
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22525 3295 22559
rect 3237 22519 3295 22525
rect 3697 22559 3755 22565
rect 3697 22525 3709 22559
rect 3743 22556 3755 22559
rect 3786 22556 3792 22568
rect 3743 22528 3792 22556
rect 3743 22525 3755 22528
rect 3697 22519 3755 22525
rect 3786 22516 3792 22528
rect 3844 22516 3850 22568
rect 4614 22516 4620 22568
rect 4672 22516 4678 22568
rect 6641 22559 6699 22565
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 6822 22556 6828 22568
rect 6687 22528 6828 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 6917 22559 6975 22565
rect 6917 22525 6929 22559
rect 6963 22556 6975 22559
rect 7168 22559 7226 22565
rect 7168 22556 7180 22559
rect 6963 22528 7180 22556
rect 6963 22525 6975 22528
rect 6917 22519 6975 22525
rect 7168 22525 7180 22528
rect 7214 22525 7226 22559
rect 7168 22519 7226 22525
rect 7653 22559 7711 22565
rect 7653 22525 7665 22559
rect 7699 22556 7711 22559
rect 7742 22556 7748 22568
rect 7699 22528 7748 22556
rect 7699 22525 7711 22528
rect 7653 22519 7711 22525
rect 7742 22516 7748 22528
rect 7800 22556 7806 22568
rect 11054 22556 11060 22568
rect 7800 22528 11060 22556
rect 7800 22516 7806 22528
rect 11054 22516 11060 22528
rect 11112 22516 11118 22568
rect 1946 22448 1952 22500
rect 2004 22488 2010 22500
rect 4632 22488 4660 22516
rect 2004 22460 4660 22488
rect 2004 22448 2010 22460
rect 8754 22448 8760 22500
rect 8812 22448 8818 22500
rect 11348 22488 11376 22587
rect 11422 22516 11428 22568
rect 11480 22556 11486 22568
rect 11793 22559 11851 22565
rect 11793 22556 11805 22559
rect 11480 22528 11805 22556
rect 11480 22516 11486 22528
rect 11793 22525 11805 22528
rect 11839 22525 11851 22559
rect 11900 22556 11928 22587
rect 11974 22584 11980 22636
rect 12032 22584 12038 22636
rect 16022 22584 16028 22636
rect 16080 22584 16086 22636
rect 16114 22584 16120 22636
rect 16172 22584 16178 22636
rect 16224 22633 16252 22664
rect 17129 22661 17141 22664
rect 17175 22661 17187 22695
rect 17129 22655 17187 22661
rect 17218 22652 17224 22704
rect 17276 22701 17282 22704
rect 17276 22695 17304 22701
rect 17292 22661 17304 22695
rect 17276 22655 17304 22661
rect 17276 22652 17282 22655
rect 17954 22652 17960 22704
rect 18012 22692 18018 22704
rect 18417 22695 18475 22701
rect 18417 22692 18429 22695
rect 18012 22664 18429 22692
rect 18012 22652 18018 22664
rect 18417 22661 18429 22664
rect 18463 22661 18475 22695
rect 18417 22655 18475 22661
rect 18598 22652 18604 22704
rect 18656 22692 18662 22704
rect 19536 22692 19564 22732
rect 18656 22664 19564 22692
rect 18656 22652 18662 22664
rect 16209 22627 16267 22633
rect 16209 22593 16221 22627
rect 16255 22593 16267 22627
rect 16209 22587 16267 22593
rect 16393 22627 16451 22633
rect 16393 22593 16405 22627
rect 16439 22624 16451 22627
rect 18322 22624 18328 22636
rect 16439 22596 16712 22624
rect 16439 22593 16451 22596
rect 16393 22587 16451 22593
rect 11900 22528 12020 22556
rect 11793 22519 11851 22525
rect 11517 22491 11575 22497
rect 11517 22488 11529 22491
rect 11348 22460 11529 22488
rect 11517 22457 11529 22460
rect 11563 22457 11575 22491
rect 11992 22488 12020 22528
rect 12066 22516 12072 22568
rect 12124 22556 12130 22568
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 12124 22528 13553 22556
rect 12124 22516 12130 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13541 22519 13599 22525
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 16224 22556 16252 22587
rect 16684 22568 16712 22596
rect 17420 22596 18328 22624
rect 15620 22528 16252 22556
rect 15620 22516 15626 22528
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16724 22528 16773 22556
rect 16724 22516 16730 22528
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 16761 22519 16819 22525
rect 12250 22488 12256 22500
rect 11992 22460 12256 22488
rect 11517 22451 11575 22457
rect 12250 22448 12256 22460
rect 12308 22448 12314 22500
rect 3602 22380 3608 22432
rect 3660 22420 3666 22432
rect 4341 22423 4399 22429
rect 4341 22420 4353 22423
rect 3660 22392 4353 22420
rect 3660 22380 3666 22392
rect 4341 22389 4353 22392
rect 4387 22389 4399 22423
rect 4341 22383 4399 22389
rect 4525 22423 4583 22429
rect 4525 22389 4537 22423
rect 4571 22420 4583 22423
rect 4614 22420 4620 22432
rect 4571 22392 4620 22420
rect 4571 22389 4583 22392
rect 4525 22383 4583 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 4890 22380 4896 22432
rect 4948 22420 4954 22432
rect 5350 22420 5356 22432
rect 4948 22392 5356 22420
rect 4948 22380 4954 22392
rect 5350 22380 5356 22392
rect 5408 22420 5414 22432
rect 5997 22423 6055 22429
rect 5997 22420 6009 22423
rect 5408 22392 6009 22420
rect 5408 22380 5414 22392
rect 5997 22389 6009 22392
rect 6043 22389 6055 22423
rect 5997 22383 6055 22389
rect 11241 22423 11299 22429
rect 11241 22389 11253 22423
rect 11287 22420 11299 22423
rect 11698 22420 11704 22432
rect 11287 22392 11704 22420
rect 11287 22389 11299 22392
rect 11241 22383 11299 22389
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 11882 22380 11888 22432
rect 11940 22380 11946 22432
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 12345 22423 12403 22429
rect 12345 22420 12357 22423
rect 12032 22392 12357 22420
rect 12032 22380 12038 22392
rect 12345 22389 12357 22392
rect 12391 22389 12403 22423
rect 12345 22383 12403 22389
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 15470 22420 15476 22432
rect 13872 22392 15476 22420
rect 13872 22380 13878 22392
rect 15470 22380 15476 22392
rect 15528 22380 15534 22432
rect 16776 22420 16804 22519
rect 17034 22516 17040 22568
rect 17092 22516 17098 22568
rect 17420 22497 17448 22596
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18509 22627 18567 22633
rect 18509 22593 18521 22627
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 17586 22516 17592 22568
rect 17644 22556 17650 22568
rect 18524 22556 18552 22587
rect 18690 22584 18696 22636
rect 18748 22584 18754 22636
rect 18966 22584 18972 22636
rect 19024 22584 19030 22636
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19245 22627 19303 22633
rect 19245 22624 19257 22627
rect 19208 22596 19257 22624
rect 19208 22584 19214 22596
rect 19245 22593 19257 22596
rect 19291 22593 19303 22627
rect 19245 22587 19303 22593
rect 19334 22584 19340 22636
rect 19392 22584 19398 22636
rect 19536 22633 19564 22664
rect 19610 22652 19616 22704
rect 19668 22692 19674 22704
rect 20180 22701 20208 22732
rect 20651 22729 20663 22763
rect 20697 22760 20709 22763
rect 20806 22760 20812 22772
rect 20697 22732 20812 22760
rect 20697 22729 20709 22732
rect 20651 22723 20709 22729
rect 20806 22720 20812 22732
rect 20864 22760 20870 22772
rect 21269 22763 21327 22769
rect 21269 22760 21281 22763
rect 20864 22732 21281 22760
rect 20864 22720 20870 22732
rect 21269 22729 21281 22732
rect 21315 22760 21327 22763
rect 21910 22760 21916 22772
rect 21315 22732 21916 22760
rect 21315 22729 21327 22732
rect 21269 22723 21327 22729
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 24765 22763 24823 22769
rect 24765 22729 24777 22763
rect 24811 22729 24823 22763
rect 24765 22723 24823 22729
rect 19705 22695 19763 22701
rect 19705 22692 19717 22695
rect 19668 22664 19717 22692
rect 19668 22652 19674 22664
rect 19705 22661 19717 22664
rect 19751 22661 19763 22695
rect 20165 22695 20223 22701
rect 19705 22655 19763 22661
rect 19935 22661 19993 22667
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22593 19579 22627
rect 19935 22627 19947 22661
rect 19981 22658 19993 22661
rect 20165 22661 20177 22695
rect 20211 22661 20223 22695
rect 19981 22627 20008 22658
rect 20165 22655 20223 22661
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 20441 22695 20499 22701
rect 20441 22692 20453 22695
rect 20404 22664 20453 22692
rect 20404 22652 20410 22664
rect 20441 22661 20453 22664
rect 20487 22661 20499 22695
rect 20441 22655 20499 22661
rect 19935 22624 20008 22627
rect 20806 22624 20812 22636
rect 19935 22621 20812 22624
rect 19980 22596 20812 22621
rect 19521 22587 19579 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 23385 22627 23443 22633
rect 23385 22593 23397 22627
rect 23431 22624 23443 22627
rect 23474 22624 23480 22636
rect 23431 22596 23480 22624
rect 23431 22593 23443 22596
rect 23385 22587 23443 22593
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 23652 22627 23710 22633
rect 23652 22593 23664 22627
rect 23698 22624 23710 22627
rect 24394 22624 24400 22636
rect 23698 22596 24400 22624
rect 23698 22593 23710 22596
rect 23652 22587 23710 22593
rect 24394 22584 24400 22596
rect 24452 22584 24458 22636
rect 24780 22624 24808 22723
rect 25222 22624 25228 22636
rect 24780 22596 25228 22624
rect 25222 22584 25228 22596
rect 25280 22624 25286 22636
rect 25409 22627 25467 22633
rect 25409 22624 25421 22627
rect 25280 22596 25421 22624
rect 25280 22584 25286 22596
rect 25409 22593 25421 22596
rect 25455 22593 25467 22627
rect 25409 22587 25467 22593
rect 25590 22584 25596 22636
rect 25648 22584 25654 22636
rect 17644 22528 18552 22556
rect 17644 22516 17650 22528
rect 17405 22491 17463 22497
rect 17405 22457 17417 22491
rect 17451 22457 17463 22491
rect 17405 22451 17463 22457
rect 17497 22491 17555 22497
rect 17497 22457 17509 22491
rect 17543 22457 17555 22491
rect 17497 22451 17555 22457
rect 17512 22420 17540 22451
rect 17678 22448 17684 22500
rect 17736 22488 17742 22500
rect 18785 22491 18843 22497
rect 18785 22488 18797 22491
rect 17736 22460 18797 22488
rect 17736 22448 17742 22460
rect 18785 22457 18797 22460
rect 18831 22457 18843 22491
rect 19352 22488 19380 22584
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 21634 22556 21640 22568
rect 19484 22528 21640 22556
rect 19484 22516 19490 22528
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 24762 22516 24768 22568
rect 24820 22556 24826 22568
rect 24857 22559 24915 22565
rect 24857 22556 24869 22559
rect 24820 22528 24869 22556
rect 24820 22516 24826 22528
rect 24857 22525 24869 22528
rect 24903 22525 24915 22559
rect 24857 22519 24915 22525
rect 18785 22451 18843 22457
rect 19076 22460 20024 22488
rect 16776 22392 17540 22420
rect 17862 22380 17868 22432
rect 17920 22380 17926 22432
rect 18049 22423 18107 22429
rect 18049 22389 18061 22423
rect 18095 22420 18107 22423
rect 19076 22420 19104 22460
rect 19996 22432 20024 22460
rect 20346 22448 20352 22500
rect 20404 22488 20410 22500
rect 20901 22491 20959 22497
rect 20901 22488 20913 22491
rect 20404 22460 20913 22488
rect 20404 22448 20410 22460
rect 20901 22457 20913 22460
rect 20947 22488 20959 22491
rect 21082 22488 21088 22500
rect 20947 22460 21088 22488
rect 20947 22457 20959 22460
rect 20901 22451 20959 22457
rect 21082 22448 21088 22460
rect 21140 22448 21146 22500
rect 18095 22392 19104 22420
rect 18095 22389 18107 22392
rect 18049 22383 18107 22389
rect 19150 22380 19156 22432
rect 19208 22380 19214 22432
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 19794 22420 19800 22432
rect 19576 22392 19800 22420
rect 19576 22380 19582 22392
rect 19794 22380 19800 22392
rect 19852 22380 19858 22432
rect 19978 22380 19984 22432
rect 20036 22380 20042 22432
rect 20625 22423 20683 22429
rect 20625 22389 20637 22423
rect 20671 22420 20683 22423
rect 20714 22420 20720 22432
rect 20671 22392 20720 22420
rect 20671 22389 20683 22392
rect 20625 22383 20683 22389
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 20809 22423 20867 22429
rect 20809 22389 20821 22423
rect 20855 22420 20867 22423
rect 20990 22420 20996 22432
rect 20855 22392 20996 22420
rect 20855 22389 20867 22392
rect 20809 22383 20867 22389
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 21174 22380 21180 22432
rect 21232 22420 21238 22432
rect 21269 22423 21327 22429
rect 21269 22420 21281 22423
rect 21232 22392 21281 22420
rect 21232 22380 21238 22392
rect 21269 22389 21281 22392
rect 21315 22420 21327 22423
rect 21358 22420 21364 22432
rect 21315 22392 21364 22420
rect 21315 22389 21327 22392
rect 21269 22383 21327 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 21450 22380 21456 22432
rect 21508 22380 21514 22432
rect 25774 22380 25780 22432
rect 25832 22380 25838 22432
rect 1104 22330 26220 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 26220 22330
rect 1104 22256 26220 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 4522 22216 4528 22228
rect 3660 22188 4528 22216
rect 3660 22176 3666 22188
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 4801 22219 4859 22225
rect 4801 22216 4813 22219
rect 4764 22188 4813 22216
rect 4764 22176 4770 22188
rect 4801 22185 4813 22188
rect 4847 22185 4859 22219
rect 4801 22179 4859 22185
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 17589 22219 17647 22225
rect 5500 22188 7604 22216
rect 5500 22176 5506 22188
rect 2774 22108 2780 22160
rect 2832 22148 2838 22160
rect 3694 22148 3700 22160
rect 2832 22120 3700 22148
rect 2832 22108 2838 22120
rect 3694 22108 3700 22120
rect 3752 22108 3758 22160
rect 3786 22108 3792 22160
rect 3844 22148 3850 22160
rect 5166 22148 5172 22160
rect 3844 22120 5172 22148
rect 3844 22108 3850 22120
rect 5166 22108 5172 22120
rect 5224 22108 5230 22160
rect 5261 22151 5319 22157
rect 5261 22117 5273 22151
rect 5307 22148 5319 22151
rect 6362 22148 6368 22160
rect 5307 22120 6368 22148
rect 5307 22117 5319 22120
rect 5261 22111 5319 22117
rect 6362 22108 6368 22120
rect 6420 22108 6426 22160
rect 7576 22148 7604 22188
rect 17589 22185 17601 22219
rect 17635 22216 17647 22219
rect 17862 22216 17868 22228
rect 17635 22188 17868 22216
rect 17635 22185 17647 22188
rect 17589 22179 17647 22185
rect 17862 22176 17868 22188
rect 17920 22176 17926 22228
rect 17957 22219 18015 22225
rect 17957 22185 17969 22219
rect 18003 22216 18015 22219
rect 18966 22216 18972 22228
rect 18003 22188 18972 22216
rect 18003 22185 18015 22188
rect 17957 22179 18015 22185
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 19334 22176 19340 22228
rect 19392 22216 19398 22228
rect 19610 22216 19616 22228
rect 19392 22188 19616 22216
rect 19392 22176 19398 22188
rect 19610 22176 19616 22188
rect 19668 22176 19674 22228
rect 20073 22219 20131 22225
rect 20073 22185 20085 22219
rect 20119 22216 20131 22219
rect 20162 22216 20168 22228
rect 20119 22188 20168 22216
rect 20119 22185 20131 22188
rect 20073 22179 20131 22185
rect 20162 22176 20168 22188
rect 20220 22216 20226 22228
rect 21358 22216 21364 22228
rect 20220 22188 20668 22216
rect 20220 22176 20226 22188
rect 8662 22148 8668 22160
rect 7576 22120 8668 22148
rect 2498 22040 2504 22092
rect 2556 22040 2562 22092
rect 2792 22080 2820 22108
rect 2608 22052 2820 22080
rect 4724 22052 5764 22080
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 2608 22012 2636 22052
rect 2464 21984 2636 22012
rect 2464 21972 2470 21984
rect 2682 21972 2688 22024
rect 2740 22012 2746 22024
rect 2777 22015 2835 22021
rect 2777 22012 2789 22015
rect 2740 21984 2789 22012
rect 2740 21972 2746 21984
rect 2777 21981 2789 21984
rect 2823 22012 2835 22015
rect 3142 22012 3148 22024
rect 2823 21984 3148 22012
rect 2823 21981 2835 21984
rect 2777 21975 2835 21981
rect 3142 21972 3148 21984
rect 3200 21972 3206 22024
rect 4614 21972 4620 22024
rect 4672 22012 4678 22024
rect 4724 22012 4752 22052
rect 4672 21984 4752 22012
rect 4801 22015 4859 22021
rect 4672 21972 4678 21984
rect 4801 21981 4813 22015
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 2292 21947 2350 21953
rect 2292 21913 2304 21947
rect 2338 21944 2350 21947
rect 3602 21944 3608 21956
rect 2338 21916 3608 21944
rect 2338 21913 2350 21916
rect 2292 21907 2350 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 2130 21836 2136 21888
rect 2188 21836 2194 21888
rect 4816 21876 4844 21975
rect 4890 21972 4896 22024
rect 4948 21972 4954 22024
rect 5074 21972 5080 22024
rect 5132 21972 5138 22024
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 5224 21984 5641 22012
rect 5224 21972 5230 21984
rect 5629 21981 5641 21984
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5092 21944 5120 21972
rect 5537 21947 5595 21953
rect 5537 21944 5549 21947
rect 5092 21916 5549 21944
rect 5537 21913 5549 21916
rect 5583 21913 5595 21947
rect 5736 21944 5764 22052
rect 5994 22040 6000 22092
rect 6052 22040 6058 22092
rect 7576 22089 7604 22120
rect 8662 22108 8668 22120
rect 8720 22108 8726 22160
rect 12250 22148 12256 22160
rect 10520 22120 12256 22148
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 6104 22052 6285 22080
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 6104 22021 6132 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 7561 22083 7619 22089
rect 7561 22080 7573 22083
rect 7539 22052 7573 22080
rect 6273 22043 6331 22049
rect 7561 22049 7573 22052
rect 7607 22049 7619 22083
rect 7561 22043 7619 22049
rect 10413 22083 10471 22089
rect 10413 22049 10425 22083
rect 10459 22080 10471 22083
rect 10520 22080 10548 22120
rect 12250 22108 12256 22120
rect 12308 22108 12314 22160
rect 16485 22151 16543 22157
rect 16485 22148 16497 22151
rect 16132 22120 16497 22148
rect 16132 22092 16160 22120
rect 16485 22117 16497 22120
rect 16531 22148 16543 22151
rect 17221 22151 17279 22157
rect 17221 22148 17233 22151
rect 16531 22120 17233 22148
rect 16531 22117 16543 22120
rect 16485 22111 16543 22117
rect 17221 22117 17233 22120
rect 17267 22117 17279 22151
rect 17221 22111 17279 22117
rect 17310 22108 17316 22160
rect 17368 22148 17374 22160
rect 18417 22151 18475 22157
rect 18417 22148 18429 22151
rect 17368 22120 18429 22148
rect 17368 22108 17374 22120
rect 18417 22117 18429 22120
rect 18463 22148 18475 22151
rect 19426 22148 19432 22160
rect 18463 22120 19432 22148
rect 18463 22117 18475 22120
rect 18417 22111 18475 22117
rect 19426 22108 19432 22120
rect 19484 22108 19490 22160
rect 20640 22157 20668 22188
rect 20916 22188 21364 22216
rect 20625 22151 20683 22157
rect 20625 22117 20637 22151
rect 20671 22117 20683 22151
rect 20625 22111 20683 22117
rect 10459 22052 10548 22080
rect 10597 22083 10655 22089
rect 10459 22049 10471 22052
rect 10413 22043 10471 22049
rect 10597 22049 10609 22083
rect 10643 22080 10655 22083
rect 10873 22083 10931 22089
rect 10873 22080 10885 22083
rect 10643 22052 10885 22080
rect 10643 22049 10655 22052
rect 10597 22043 10655 22049
rect 10873 22049 10885 22052
rect 10919 22049 10931 22083
rect 10873 22043 10931 22049
rect 11146 22040 11152 22092
rect 11204 22080 11210 22092
rect 11204 22052 11836 22080
rect 11204 22040 11210 22052
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 6196 21944 6224 21975
rect 6362 21972 6368 22024
rect 6420 21972 6426 22024
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 8297 22015 8355 22021
rect 8297 22012 8309 22015
rect 7156 21984 8309 22012
rect 7156 21972 7162 21984
rect 8297 21981 8309 21984
rect 8343 21981 8355 22015
rect 8297 21975 8355 21981
rect 8481 22015 8539 22021
rect 8481 21981 8493 22015
rect 8527 22012 8539 22015
rect 9122 22012 9128 22024
rect 8527 21984 9128 22012
rect 8527 21981 8539 21984
rect 8481 21975 8539 21981
rect 9122 21972 9128 21984
rect 9180 21972 9186 22024
rect 10505 22015 10563 22021
rect 10505 21981 10517 22015
rect 10551 21981 10563 22015
rect 10505 21975 10563 21981
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 5736 21916 6224 21944
rect 8046 21947 8104 21953
rect 5537 21907 5595 21913
rect 8046 21913 8058 21947
rect 8092 21944 8104 21947
rect 8389 21947 8447 21953
rect 8389 21944 8401 21947
rect 8092 21916 8401 21944
rect 8092 21913 8104 21916
rect 8046 21907 8104 21913
rect 8389 21913 8401 21916
rect 8435 21913 8447 21947
rect 8389 21907 8447 21913
rect 4991 21879 5049 21885
rect 4991 21876 5003 21879
rect 4816 21848 5003 21876
rect 4991 21845 5003 21848
rect 5037 21845 5049 21879
rect 4991 21839 5049 21845
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 5408 21848 5457 21876
rect 5408 21836 5414 21848
rect 5445 21845 5457 21848
rect 5491 21845 5503 21879
rect 5445 21839 5503 21845
rect 5813 21879 5871 21885
rect 5813 21845 5825 21879
rect 5859 21876 5871 21879
rect 5902 21876 5908 21888
rect 5859 21848 5908 21876
rect 5859 21845 5871 21848
rect 5813 21839 5871 21845
rect 5902 21836 5908 21848
rect 5960 21876 5966 21888
rect 6822 21876 6828 21888
rect 5960 21848 6828 21876
rect 5960 21836 5966 21848
rect 6822 21836 6828 21848
rect 6880 21836 6886 21888
rect 7834 21836 7840 21888
rect 7892 21836 7898 21888
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 8202 21836 8208 21888
rect 8260 21836 8266 21888
rect 10134 21836 10140 21888
rect 10192 21876 10198 21888
rect 10229 21879 10287 21885
rect 10229 21876 10241 21879
rect 10192 21848 10241 21876
rect 10192 21836 10198 21848
rect 10229 21845 10241 21848
rect 10275 21845 10287 21879
rect 10520 21876 10548 21975
rect 10704 21944 10732 21975
rect 11238 21972 11244 22024
rect 11296 22012 11302 22024
rect 11422 22012 11428 22024
rect 11296 21984 11428 22012
rect 11296 21972 11302 21984
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 11698 21944 11704 21956
rect 10704 21916 11704 21944
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 11808 21944 11836 22052
rect 12176 22052 12572 22080
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 12176 22021 12204 22052
rect 12544 22024 12572 22052
rect 16114 22040 16120 22092
rect 16172 22040 16178 22092
rect 16666 22040 16672 22092
rect 16724 22080 16730 22092
rect 16945 22083 17003 22089
rect 16945 22080 16957 22083
rect 16724 22052 16957 22080
rect 16724 22040 16730 22052
rect 16945 22049 16957 22052
rect 16991 22049 17003 22083
rect 18046 22080 18052 22092
rect 16945 22043 17003 22049
rect 17696 22052 18052 22080
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11940 21984 12173 22012
rect 11940 21972 11946 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 12342 21972 12348 22024
rect 12400 21972 12406 22024
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12437 21947 12495 21953
rect 12437 21944 12449 21947
rect 11808 21916 12449 21944
rect 12437 21913 12449 21916
rect 12483 21944 12495 21947
rect 12636 21944 12664 21975
rect 12802 21972 12808 22024
rect 12860 21972 12866 22024
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13596 21984 14105 22012
rect 13596 21972 13602 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 16025 22015 16083 22021
rect 16025 22012 16037 22015
rect 15620 21984 16037 22012
rect 15620 21972 15626 21984
rect 16025 21981 16037 21984
rect 16071 21981 16083 22015
rect 16132 22012 16160 22040
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 16132 21984 16221 22012
rect 16025 21975 16083 21981
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 16301 22015 16359 22021
rect 16301 21981 16313 22015
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16485 22015 16543 22021
rect 16485 21981 16497 22015
rect 16531 22012 16543 22015
rect 17034 22012 17040 22024
rect 16531 21984 17040 22012
rect 16531 21981 16543 21984
rect 16485 21975 16543 21981
rect 12483 21916 12664 21944
rect 16316 21944 16344 21975
rect 17034 21972 17040 21984
rect 17092 22012 17098 22024
rect 17092 21984 17172 22012
rect 17092 21972 17098 21984
rect 16758 21944 16764 21956
rect 16316 21916 16764 21944
rect 12483 21913 12495 21916
rect 12437 21907 12495 21913
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 17144 21944 17172 21984
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 17586 22012 17592 22024
rect 17276 21984 17592 22012
rect 17276 21972 17282 21984
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 17696 22021 17724 22052
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 20346 22080 20352 22092
rect 20072 22052 20352 22080
rect 17681 22015 17739 22021
rect 17681 21981 17693 22015
rect 17727 21981 17739 22015
rect 17681 21975 17739 21981
rect 17865 22015 17923 22021
rect 17865 21981 17877 22015
rect 17911 21981 17923 22015
rect 17865 21975 17923 21981
rect 18692 22015 18750 22021
rect 18692 21981 18704 22015
rect 18738 21981 18750 22015
rect 18692 21975 18750 21981
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 22012 18843 22015
rect 19058 22012 19064 22024
rect 18831 21984 19064 22012
rect 18831 21981 18843 21984
rect 18785 21975 18843 21981
rect 17880 21944 17908 21975
rect 17144 21916 17908 21944
rect 18708 21944 18736 21975
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 20072 21987 20100 22052
rect 20346 22040 20352 22052
rect 20404 22040 20410 22092
rect 20640 22080 20668 22111
rect 20714 22108 20720 22160
rect 20772 22148 20778 22160
rect 20916 22148 20944 22188
rect 21358 22176 21364 22188
rect 21416 22176 21422 22228
rect 21542 22176 21548 22228
rect 21600 22216 21606 22228
rect 21910 22216 21916 22228
rect 21600 22188 21916 22216
rect 21600 22176 21606 22188
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 22465 22219 22523 22225
rect 22465 22185 22477 22219
rect 22511 22185 22523 22219
rect 22465 22179 22523 22185
rect 20772 22120 20944 22148
rect 21085 22151 21143 22157
rect 20772 22108 20778 22120
rect 21085 22117 21097 22151
rect 21131 22148 21143 22151
rect 21174 22148 21180 22160
rect 21131 22120 21180 22148
rect 21131 22117 21143 22120
rect 21085 22111 21143 22117
rect 21174 22108 21180 22120
rect 21232 22108 21238 22160
rect 21376 22148 21404 22176
rect 22005 22151 22063 22157
rect 22005 22148 22017 22151
rect 21376 22120 22017 22148
rect 22005 22117 22017 22120
rect 22051 22117 22063 22151
rect 22005 22111 22063 22117
rect 21266 22080 21272 22092
rect 20640 22052 21272 22080
rect 21266 22040 21272 22052
rect 21324 22080 21330 22092
rect 21361 22083 21419 22089
rect 21361 22080 21373 22083
rect 21324 22052 21373 22080
rect 21324 22040 21330 22052
rect 21361 22049 21373 22052
rect 21407 22049 21419 22083
rect 21361 22043 21419 22049
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 22094 22080 22100 22092
rect 21591 22052 22100 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 22094 22040 22100 22052
rect 22152 22040 22158 22092
rect 22189 22083 22247 22089
rect 22189 22049 22201 22083
rect 22235 22080 22247 22083
rect 22480 22080 22508 22179
rect 24394 22176 24400 22228
rect 24452 22176 24458 22228
rect 22738 22080 22744 22092
rect 22235 22052 22744 22080
rect 22235 22049 22247 22052
rect 22189 22043 22247 22049
rect 22738 22040 22744 22052
rect 22796 22040 22802 22092
rect 23474 22040 23480 22092
rect 23532 22080 23538 22092
rect 24949 22083 25007 22089
rect 24949 22080 24961 22083
rect 23532 22052 24961 22080
rect 23532 22040 23538 22052
rect 24949 22049 24961 22052
rect 24995 22049 25007 22083
rect 24949 22043 25007 22049
rect 20622 22012 20628 22024
rect 20027 21981 20100 21987
rect 19702 21944 19708 21956
rect 18708 21916 19708 21944
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 20027 21947 20039 21981
rect 20073 21950 20100 21981
rect 20272 21984 20628 22012
rect 20272 21953 20300 21984
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20806 21972 20812 22024
rect 20864 22012 20870 22024
rect 21453 22015 21511 22021
rect 20864 21984 21404 22012
rect 20864 21972 20870 21984
rect 20073 21947 20085 21950
rect 20027 21941 20085 21947
rect 20257 21947 20315 21953
rect 20257 21913 20269 21947
rect 20303 21913 20315 21947
rect 20257 21907 20315 21913
rect 11146 21876 11152 21888
rect 10520 21848 11152 21876
rect 10229 21839 10287 21845
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11882 21876 11888 21888
rect 11655 21848 11888 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11882 21836 11888 21848
rect 11940 21836 11946 21888
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21876 12771 21879
rect 13170 21876 13176 21888
rect 12759 21848 13176 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 14458 21836 14464 21888
rect 14516 21876 14522 21888
rect 14642 21876 14648 21888
rect 14516 21848 14648 21876
rect 14516 21836 14522 21848
rect 14642 21836 14648 21848
rect 14700 21876 14706 21888
rect 14737 21879 14795 21885
rect 14737 21876 14749 21879
rect 14700 21848 14749 21876
rect 14700 21836 14706 21848
rect 14737 21845 14749 21848
rect 14783 21845 14795 21879
rect 14737 21839 14795 21845
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 17218 21876 17224 21888
rect 16163 21848 17224 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 17218 21836 17224 21848
rect 17276 21836 17282 21888
rect 17405 21879 17463 21885
rect 17405 21845 17417 21879
rect 17451 21876 17463 21879
rect 19794 21876 19800 21888
rect 17451 21848 19800 21876
rect 17451 21845 17463 21848
rect 17405 21839 17463 21845
rect 19794 21836 19800 21848
rect 19852 21836 19858 21888
rect 19886 21836 19892 21888
rect 19944 21836 19950 21888
rect 20806 21836 20812 21888
rect 20864 21836 20870 21888
rect 20916 21885 20944 21984
rect 21376 21956 21404 21984
rect 21453 21981 21465 22015
rect 21499 22006 21511 22015
rect 21913 22015 21971 22021
rect 21499 22002 21588 22006
rect 21499 21981 21548 22002
rect 21453 21978 21548 21981
rect 21453 21975 21511 21978
rect 21358 21904 21364 21956
rect 21416 21904 21422 21956
rect 21542 21950 21548 21978
rect 21600 21950 21606 22002
rect 21913 21981 21925 22015
rect 21959 21981 21971 22015
rect 22112 22012 22140 22040
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22112 21984 22293 22012
rect 21913 21975 21971 21981
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 21928 21944 21956 21975
rect 24762 21972 24768 22024
rect 24820 21972 24826 22024
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 21652 21916 21956 21944
rect 20901 21879 20959 21885
rect 20901 21845 20913 21879
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 21652 21876 21680 21916
rect 23658 21904 23664 21956
rect 23716 21944 23722 21956
rect 25240 21944 25268 21975
rect 25590 21972 25596 22024
rect 25648 21972 25654 22024
rect 23716 21916 25268 21944
rect 23716 21904 23722 21916
rect 21232 21848 21680 21876
rect 21821 21879 21879 21885
rect 21232 21836 21238 21848
rect 21821 21845 21833 21879
rect 21867 21876 21879 21879
rect 22002 21876 22008 21888
rect 21867 21848 22008 21876
rect 21867 21845 21879 21848
rect 21821 21839 21879 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22189 21879 22247 21885
rect 22189 21845 22201 21879
rect 22235 21876 22247 21879
rect 22370 21876 22376 21888
rect 22235 21848 22376 21876
rect 22235 21845 22247 21848
rect 22189 21839 22247 21845
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 23934 21836 23940 21888
rect 23992 21876 23998 21888
rect 24857 21879 24915 21885
rect 24857 21876 24869 21879
rect 23992 21848 24869 21876
rect 23992 21836 23998 21848
rect 24857 21845 24869 21848
rect 24903 21845 24915 21879
rect 24857 21839 24915 21845
rect 25406 21836 25412 21888
rect 25464 21836 25470 21888
rect 25777 21879 25835 21885
rect 25777 21845 25789 21879
rect 25823 21876 25835 21879
rect 25958 21876 25964 21888
rect 25823 21848 25964 21876
rect 25823 21845 25835 21848
rect 25777 21839 25835 21845
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 1104 21786 26220 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 26220 21786
rect 1104 21712 26220 21734
rect 3602 21632 3608 21684
rect 3660 21632 3666 21684
rect 6914 21672 6920 21684
rect 6840 21644 6920 21672
rect 2130 21564 2136 21616
rect 2188 21604 2194 21616
rect 2286 21607 2344 21613
rect 2286 21604 2298 21607
rect 2188 21576 2298 21604
rect 2188 21564 2194 21576
rect 2286 21573 2298 21576
rect 2332 21573 2344 21607
rect 2286 21567 2344 21573
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 900 21508 1409 21536
rect 900 21496 906 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 3326 21496 3332 21548
rect 3384 21536 3390 21548
rect 3513 21539 3571 21545
rect 3513 21536 3525 21539
rect 3384 21508 3525 21536
rect 3384 21496 3390 21508
rect 3513 21505 3525 21508
rect 3559 21505 3571 21539
rect 3513 21499 3571 21505
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21536 3755 21539
rect 3786 21536 3792 21548
rect 3743 21508 3792 21536
rect 3743 21505 3755 21508
rect 3697 21499 3755 21505
rect 3786 21496 3792 21508
rect 3844 21496 3850 21548
rect 6840 21545 6868 21644
rect 6914 21632 6920 21644
rect 6972 21672 6978 21684
rect 7393 21675 7451 21681
rect 7393 21672 7405 21675
rect 6972 21644 7405 21672
rect 6972 21632 6978 21644
rect 7393 21641 7405 21644
rect 7439 21641 7451 21675
rect 7393 21635 7451 21641
rect 7561 21675 7619 21681
rect 7561 21641 7573 21675
rect 7607 21672 7619 21675
rect 9122 21672 9128 21684
rect 7607 21644 9128 21672
rect 7607 21641 7619 21644
rect 7561 21635 7619 21641
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 11333 21675 11391 21681
rect 11333 21641 11345 21675
rect 11379 21672 11391 21675
rect 11790 21672 11796 21684
rect 11379 21644 11796 21672
rect 11379 21641 11391 21644
rect 11333 21635 11391 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12250 21632 12256 21684
rect 12308 21672 12314 21684
rect 12802 21672 12808 21684
rect 12308 21644 12808 21672
rect 12308 21632 12314 21644
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 13538 21632 13544 21684
rect 13596 21632 13602 21684
rect 22186 21672 22192 21684
rect 20456 21644 22192 21672
rect 7193 21607 7251 21613
rect 7193 21573 7205 21607
rect 7239 21573 7251 21607
rect 8294 21604 8300 21616
rect 7193 21567 7251 21573
rect 7668 21576 8300 21604
rect 6825 21539 6883 21545
rect 6825 21505 6837 21539
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21505 6975 21539
rect 6917 21499 6975 21505
rect 1946 21428 1952 21480
rect 2004 21468 2010 21480
rect 2041 21471 2099 21477
rect 2041 21468 2053 21471
rect 2004 21440 2053 21468
rect 2004 21428 2010 21440
rect 2041 21437 2053 21440
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 6840 21468 6868 21499
rect 6788 21440 6868 21468
rect 6788 21428 6794 21440
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 3234 21332 3240 21344
rect 1627 21304 3240 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 3418 21292 3424 21344
rect 3476 21292 3482 21344
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 6638 21332 6644 21344
rect 6512 21304 6644 21332
rect 6512 21292 6518 21304
rect 6638 21292 6644 21304
rect 6696 21332 6702 21344
rect 6932 21332 6960 21499
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 7101 21539 7159 21545
rect 7101 21536 7113 21539
rect 7064 21508 7113 21536
rect 7064 21496 7070 21508
rect 7101 21505 7113 21508
rect 7147 21536 7159 21539
rect 7208 21536 7236 21567
rect 7668 21545 7696 21576
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 12710 21564 12716 21616
rect 12768 21604 12774 21616
rect 13446 21604 13452 21616
rect 12768 21576 13452 21604
rect 12768 21564 12774 21576
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 7147 21508 7236 21536
rect 7147 21505 7159 21508
rect 7101 21499 7159 21505
rect 7098 21360 7104 21412
rect 7156 21360 7162 21412
rect 7208 21400 7236 21508
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 7920 21539 7978 21545
rect 7920 21505 7932 21539
rect 7966 21536 7978 21539
rect 8202 21536 8208 21548
rect 7966 21508 8208 21536
rect 7966 21505 7978 21508
rect 7920 21499 7978 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 10220 21539 10278 21545
rect 10220 21505 10232 21539
rect 10266 21536 10278 21539
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 10266 21508 11529 21536
rect 10266 21505 10278 21508
rect 10220 21499 10278 21505
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11974 21496 11980 21548
rect 12032 21496 12038 21548
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12336 21539 12394 21545
rect 12336 21505 12348 21539
rect 12382 21536 12394 21539
rect 12894 21536 12900 21548
rect 12382 21508 12900 21536
rect 12382 21505 12394 21508
rect 12336 21499 12394 21505
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 9582 21428 9588 21480
rect 9640 21468 9646 21480
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9640 21440 9965 21468
rect 9640 21428 9646 21440
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 9953 21431 10011 21437
rect 13556 21400 13584 21632
rect 20349 21607 20407 21613
rect 20349 21604 20361 21607
rect 7208 21372 7696 21400
rect 7377 21335 7435 21341
rect 7377 21332 7389 21335
rect 6696 21304 7389 21332
rect 6696 21292 6702 21304
rect 7377 21301 7389 21304
rect 7423 21301 7435 21335
rect 7668 21332 7696 21372
rect 13372 21372 13584 21400
rect 13648 21576 15792 21604
rect 9033 21335 9091 21341
rect 9033 21332 9045 21335
rect 7668 21304 9045 21332
rect 7377 21295 7435 21301
rect 9033 21301 9045 21304
rect 9079 21332 9091 21335
rect 9490 21332 9496 21344
rect 9079 21304 9496 21332
rect 9079 21301 9091 21304
rect 9033 21295 9091 21301
rect 9490 21292 9496 21304
rect 9548 21292 9554 21344
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 13372 21332 13400 21372
rect 13648 21344 13676 21576
rect 14665 21539 14723 21545
rect 14665 21505 14677 21539
rect 14711 21536 14723 21539
rect 14826 21536 14832 21548
rect 14711 21508 14832 21536
rect 14711 21505 14723 21508
rect 14665 21499 14723 21505
rect 14826 21496 14832 21508
rect 14884 21496 14890 21548
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21536 14979 21539
rect 15654 21536 15660 21548
rect 14967 21508 15660 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 15764 21468 15792 21576
rect 19996 21576 20361 21604
rect 19996 21548 20024 21576
rect 20349 21573 20361 21576
rect 20395 21573 20407 21607
rect 20349 21567 20407 21573
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21536 19855 21539
rect 19978 21536 19984 21548
rect 19843 21508 19984 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20456 21536 20484 21644
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 23382 21672 23388 21684
rect 22511 21644 23388 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 23492 21644 25145 21672
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21545 21607 21603 21613
rect 21545 21604 21557 21607
rect 21048 21576 21557 21604
rect 21048 21564 21054 21576
rect 21545 21573 21557 21576
rect 21591 21604 21603 21607
rect 22278 21604 22284 21616
rect 21591 21576 22284 21604
rect 21591 21573 21603 21576
rect 21545 21567 21603 21573
rect 22278 21564 22284 21576
rect 22336 21604 22342 21616
rect 22336 21576 22600 21604
rect 22336 21564 22342 21576
rect 20119 21508 20484 21536
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21536 20867 21539
rect 21174 21536 21180 21548
rect 20855 21508 21180 21536
rect 20855 21505 20867 21508
rect 20809 21499 20867 21505
rect 21174 21496 21180 21508
rect 21232 21496 21238 21548
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 21361 21539 21419 21545
rect 21361 21536 21373 21539
rect 21324 21508 21373 21536
rect 21324 21496 21330 21508
rect 21361 21505 21373 21508
rect 21407 21536 21419 21539
rect 21726 21536 21732 21548
rect 21407 21508 21732 21536
rect 21407 21505 21419 21508
rect 21361 21499 21419 21505
rect 21726 21496 21732 21508
rect 21784 21496 21790 21548
rect 21821 21539 21879 21545
rect 21821 21505 21833 21539
rect 21867 21536 21879 21539
rect 21910 21536 21916 21548
rect 21867 21508 21916 21536
rect 21867 21505 21879 21508
rect 21821 21499 21879 21505
rect 21910 21496 21916 21508
rect 21968 21496 21974 21548
rect 22002 21496 22008 21548
rect 22060 21496 22066 21548
rect 22572 21545 22600 21576
rect 22097 21539 22155 21545
rect 22097 21505 22109 21539
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 23198 21536 23204 21548
rect 22879 21508 23204 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 15611 21440 15792 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 19886 21428 19892 21480
rect 19944 21468 19950 21480
rect 20346 21468 20352 21480
rect 19944 21440 20352 21468
rect 19944 21428 19950 21440
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20714 21428 20720 21480
rect 20772 21468 20778 21480
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 20772 21440 20913 21468
rect 20772 21428 20778 21440
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 21085 21471 21143 21477
rect 21085 21437 21097 21471
rect 21131 21468 21143 21471
rect 21131 21440 21312 21468
rect 21131 21437 21143 21440
rect 21085 21431 21143 21437
rect 19978 21360 19984 21412
rect 20036 21360 20042 21412
rect 21174 21400 21180 21412
rect 20088 21372 21180 21400
rect 12308 21304 13400 21332
rect 13449 21335 13507 21341
rect 12308 21292 12314 21304
rect 13449 21301 13461 21335
rect 13495 21332 13507 21335
rect 13630 21332 13636 21344
rect 13495 21304 13636 21332
rect 13495 21301 13507 21304
rect 13449 21295 13507 21301
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 15013 21335 15071 21341
rect 15013 21332 15025 21335
rect 13872 21304 15025 21332
rect 13872 21292 13878 21304
rect 15013 21301 15025 21304
rect 15059 21301 15071 21335
rect 15013 21295 15071 21301
rect 19150 21292 19156 21344
rect 19208 21332 19214 21344
rect 20088 21332 20116 21372
rect 21174 21360 21180 21372
rect 21232 21360 21238 21412
rect 21284 21400 21312 21440
rect 21634 21428 21640 21480
rect 21692 21468 21698 21480
rect 22112 21468 22140 21499
rect 21692 21440 22140 21468
rect 21692 21428 21698 21440
rect 21284 21372 21588 21400
rect 19208 21304 20116 21332
rect 19208 21292 19214 21304
rect 20162 21292 20168 21344
rect 20220 21332 20226 21344
rect 20257 21335 20315 21341
rect 20257 21332 20269 21335
rect 20220 21304 20269 21332
rect 20220 21292 20226 21304
rect 20257 21301 20269 21304
rect 20303 21301 20315 21335
rect 20257 21295 20315 21301
rect 20625 21335 20683 21341
rect 20625 21301 20637 21335
rect 20671 21332 20683 21335
rect 20806 21332 20812 21344
rect 20671 21304 20812 21332
rect 20671 21301 20683 21304
rect 20625 21295 20683 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 20993 21335 21051 21341
rect 20993 21301 21005 21335
rect 21039 21332 21051 21335
rect 21082 21332 21088 21344
rect 21039 21304 21088 21332
rect 21039 21301 21051 21304
rect 20993 21295 21051 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 21266 21292 21272 21344
rect 21324 21292 21330 21344
rect 21560 21332 21588 21372
rect 21818 21360 21824 21412
rect 21876 21400 21882 21412
rect 22204 21400 22232 21499
rect 23198 21496 23204 21508
rect 23256 21496 23262 21548
rect 23492 21545 23520 21644
rect 25133 21641 25145 21644
rect 25179 21641 25191 21675
rect 25133 21635 25191 21641
rect 23477 21539 23535 21545
rect 23477 21505 23489 21539
rect 23523 21505 23535 21539
rect 23477 21499 23535 21505
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 23750 21536 23756 21548
rect 23624 21508 23756 21536
rect 23624 21496 23630 21508
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 24026 21545 24032 21548
rect 24020 21499 24032 21545
rect 24026 21496 24032 21499
rect 24084 21496 24090 21548
rect 25148 21536 25176 21635
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25148 21508 25789 21536
rect 25777 21505 25789 21508
rect 25823 21505 25835 21539
rect 25777 21499 25835 21505
rect 22922 21428 22928 21480
rect 22980 21428 22986 21480
rect 21876 21372 22232 21400
rect 21876 21360 21882 21372
rect 23658 21360 23664 21412
rect 23716 21360 23722 21412
rect 22554 21332 22560 21344
rect 21560 21304 22560 21332
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 25222 21292 25228 21344
rect 25280 21292 25286 21344
rect 1104 21242 26220 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 26220 21242
rect 1104 21168 26220 21190
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5350 21128 5356 21140
rect 5215 21100 5356 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 3234 20952 3240 21004
rect 3292 20992 3298 21004
rect 5184 20992 5212 21091
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 11238 21088 11244 21140
rect 11296 21088 11302 21140
rect 11974 21088 11980 21140
rect 12032 21128 12038 21140
rect 12710 21128 12716 21140
rect 12032 21100 12716 21128
rect 12032 21088 12038 21100
rect 12710 21088 12716 21100
rect 12768 21088 12774 21140
rect 12802 21088 12808 21140
rect 12860 21128 12866 21140
rect 13357 21131 13415 21137
rect 13357 21128 13369 21131
rect 12860 21100 13369 21128
rect 12860 21088 12866 21100
rect 13357 21097 13369 21100
rect 13403 21097 13415 21131
rect 13357 21091 13415 21097
rect 13446 21088 13452 21140
rect 13504 21128 13510 21140
rect 13541 21131 13599 21137
rect 13541 21128 13553 21131
rect 13504 21100 13553 21128
rect 13504 21088 13510 21100
rect 13541 21097 13553 21100
rect 13587 21128 13599 21131
rect 14090 21128 14096 21140
rect 13587 21100 14096 21128
rect 13587 21097 13599 21100
rect 13541 21091 13599 21097
rect 14090 21088 14096 21100
rect 14148 21088 14154 21140
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 14921 21131 14979 21137
rect 14921 21128 14933 21131
rect 14884 21100 14933 21128
rect 14884 21088 14890 21100
rect 14921 21097 14933 21100
rect 14967 21097 14979 21131
rect 14921 21091 14979 21097
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20349 21131 20407 21137
rect 20349 21128 20361 21131
rect 20036 21100 20361 21128
rect 20036 21088 20042 21100
rect 5537 21063 5595 21069
rect 5537 21029 5549 21063
rect 5583 21060 5595 21063
rect 5718 21060 5724 21072
rect 5583 21032 5724 21060
rect 5583 21029 5595 21032
rect 5537 21023 5595 21029
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 5810 21020 5816 21072
rect 5868 21060 5874 21072
rect 6638 21060 6644 21072
rect 5868 21032 6644 21060
rect 5868 21020 5874 21032
rect 6638 21020 6644 21032
rect 6696 21060 6702 21072
rect 6696 21032 7328 21060
rect 6696 21020 6702 21032
rect 6089 20995 6147 21001
rect 6089 20992 6101 20995
rect 3292 20964 4292 20992
rect 3292 20952 3298 20964
rect 1857 20927 1915 20933
rect 1857 20893 1869 20927
rect 1903 20924 1915 20927
rect 1946 20924 1952 20936
rect 1903 20896 1952 20924
rect 1903 20893 1915 20896
rect 1857 20887 1915 20893
rect 1946 20884 1952 20896
rect 2004 20924 2010 20936
rect 2406 20924 2412 20936
rect 2004 20896 2412 20924
rect 2004 20884 2010 20896
rect 2406 20884 2412 20896
rect 2464 20884 2470 20936
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 3329 20927 3387 20933
rect 3329 20924 3341 20927
rect 2924 20896 3341 20924
rect 2924 20884 2930 20896
rect 3329 20893 3341 20896
rect 3375 20893 3387 20927
rect 3329 20887 3387 20893
rect 3418 20884 3424 20936
rect 3476 20924 3482 20936
rect 3513 20927 3571 20933
rect 3513 20924 3525 20927
rect 3476 20896 3525 20924
rect 3476 20884 3482 20896
rect 3513 20893 3525 20896
rect 3559 20924 3571 20927
rect 4062 20924 4068 20936
rect 3559 20896 4068 20924
rect 3559 20893 3571 20896
rect 3513 20887 3571 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4264 20933 4292 20964
rect 5000 20964 5212 20992
rect 5368 20964 6101 20992
rect 5000 20933 5028 20964
rect 5368 20933 5396 20964
rect 6089 20961 6101 20964
rect 6135 20992 6147 20995
rect 6362 20992 6368 21004
rect 6135 20964 6368 20992
rect 6135 20961 6147 20964
rect 6089 20955 6147 20961
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 6454 20952 6460 21004
rect 6512 20992 6518 21004
rect 7193 20995 7251 21001
rect 7193 20992 7205 20995
rect 6512 20964 7205 20992
rect 6512 20952 6518 20964
rect 7193 20961 7205 20964
rect 7239 20961 7251 20995
rect 7193 20955 7251 20961
rect 4249 20927 4307 20933
rect 4249 20893 4261 20927
rect 4295 20893 4307 20927
rect 4249 20887 4307 20893
rect 4892 20927 4950 20933
rect 4892 20893 4904 20927
rect 4938 20893 4950 20927
rect 4892 20887 4950 20893
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 5077 20927 5135 20933
rect 5077 20893 5089 20927
rect 5123 20893 5135 20927
rect 5077 20887 5135 20893
rect 5353 20927 5411 20933
rect 5353 20893 5365 20927
rect 5399 20893 5411 20927
rect 5353 20887 5411 20893
rect 2130 20865 2136 20868
rect 2124 20819 2136 20865
rect 2130 20816 2136 20819
rect 2188 20816 2194 20868
rect 4798 20856 4804 20868
rect 4448 20828 4804 20856
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 4448 20797 4476 20828
rect 4798 20816 4804 20828
rect 4856 20856 4862 20868
rect 4899 20856 4927 20887
rect 5092 20856 5120 20887
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20924 5963 20927
rect 5994 20924 6000 20936
rect 5951 20896 6000 20924
rect 5951 20893 5963 20896
rect 5905 20887 5963 20893
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6181 20927 6239 20933
rect 6181 20893 6193 20927
rect 6227 20924 6239 20927
rect 6273 20927 6331 20933
rect 6273 20924 6285 20927
rect 6227 20896 6285 20924
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6273 20893 6285 20896
rect 6319 20924 6331 20927
rect 6546 20924 6552 20936
rect 6319 20896 6552 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20924 7067 20927
rect 7300 20924 7328 21032
rect 9490 21020 9496 21072
rect 9548 21020 9554 21072
rect 12176 21032 12572 21060
rect 12176 20992 12204 21032
rect 11348 20964 12204 20992
rect 12544 20992 12572 21032
rect 12618 21020 12624 21072
rect 12676 21020 12682 21072
rect 14366 21020 14372 21072
rect 14424 21060 14430 21072
rect 20073 21063 20131 21069
rect 20073 21060 20085 21063
rect 14424 21032 15240 21060
rect 14424 21020 14430 21032
rect 12710 20992 12716 21004
rect 12544 20964 12716 20992
rect 8757 20927 8815 20933
rect 8757 20924 8769 20927
rect 7055 20896 7328 20924
rect 8312 20896 8769 20924
rect 7055 20893 7067 20896
rect 7009 20887 7067 20893
rect 8312 20868 8340 20896
rect 8757 20893 8769 20896
rect 8803 20924 8815 20927
rect 9582 20924 9588 20936
rect 8803 20896 9588 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 9582 20884 9588 20896
rect 9640 20924 9646 20936
rect 10134 20933 10140 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9640 20896 9873 20924
rect 9640 20884 9646 20896
rect 9861 20893 9873 20896
rect 9907 20893 9919 20927
rect 10128 20924 10140 20933
rect 10095 20896 10140 20924
rect 9861 20887 9919 20893
rect 10128 20887 10140 20896
rect 10134 20884 10140 20887
rect 10192 20884 10198 20936
rect 11348 20933 11376 20964
rect 12710 20952 12716 20964
rect 12768 20992 12774 21004
rect 12897 20995 12955 21001
rect 12897 20992 12909 20995
rect 12768 20964 12909 20992
rect 12768 20952 12774 20964
rect 12897 20961 12909 20964
rect 12943 20961 12955 20995
rect 12897 20955 12955 20961
rect 12986 20952 12992 21004
rect 13044 20952 13050 21004
rect 13081 20995 13139 21001
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13446 20992 13452 21004
rect 13127 20964 13452 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 13630 20952 13636 21004
rect 13688 20952 13694 21004
rect 14274 20952 14280 21004
rect 14332 20952 14338 21004
rect 14458 20952 14464 21004
rect 14516 20952 14522 21004
rect 15105 20995 15163 21001
rect 15105 20992 15117 20995
rect 14568 20964 15117 20992
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 11517 20927 11575 20933
rect 11517 20893 11529 20927
rect 11563 20924 11575 20927
rect 12158 20924 12164 20936
rect 11563 20896 12164 20924
rect 11563 20893 11575 20896
rect 11517 20887 11575 20893
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 12434 20884 12440 20936
rect 12492 20884 12498 20936
rect 12802 20884 12808 20936
rect 12860 20884 12866 20936
rect 13256 20927 13314 20933
rect 13256 20924 13268 20927
rect 13188 20896 13268 20924
rect 6641 20859 6699 20865
rect 6641 20856 6653 20859
rect 4856 20828 6653 20856
rect 4856 20816 4862 20828
rect 6641 20825 6653 20828
rect 6687 20825 6699 20859
rect 6641 20819 6699 20825
rect 6730 20816 6736 20868
rect 6788 20856 6794 20868
rect 6788 20828 7512 20856
rect 6788 20816 6794 20828
rect 4433 20791 4491 20797
rect 4433 20757 4445 20791
rect 4479 20757 4491 20791
rect 4433 20751 4491 20757
rect 4614 20748 4620 20800
rect 4672 20748 4678 20800
rect 5626 20748 5632 20800
rect 5684 20748 5690 20800
rect 6822 20748 6828 20800
rect 6880 20748 6886 20800
rect 7374 20748 7380 20800
rect 7432 20748 7438 20800
rect 7484 20788 7512 20828
rect 8294 20816 8300 20868
rect 8352 20816 8358 20868
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 8490 20859 8548 20865
rect 8490 20856 8502 20859
rect 8444 20828 8502 20856
rect 8444 20816 8450 20828
rect 8490 20825 8502 20828
rect 8536 20825 8548 20859
rect 8490 20819 8548 20825
rect 8938 20816 8944 20868
rect 8996 20816 9002 20868
rect 9030 20816 9036 20868
rect 9088 20856 9094 20868
rect 9217 20859 9275 20865
rect 9217 20856 9229 20859
rect 9088 20828 9229 20856
rect 9088 20816 9094 20828
rect 9217 20825 9229 20828
rect 9263 20825 9275 20859
rect 9217 20819 9275 20825
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 7484 20760 9137 20788
rect 9125 20757 9137 20760
rect 9171 20757 9183 20791
rect 9125 20751 9183 20757
rect 9306 20748 9312 20800
rect 9364 20748 9370 20800
rect 11514 20748 11520 20800
rect 11572 20748 11578 20800
rect 11882 20748 11888 20800
rect 11940 20748 11946 20800
rect 12176 20788 12204 20884
rect 13188 20788 13216 20896
rect 13256 20893 13268 20896
rect 13302 20893 13314 20927
rect 13256 20887 13314 20893
rect 13722 20884 13728 20936
rect 13780 20924 13786 20936
rect 13909 20927 13967 20933
rect 13909 20924 13921 20927
rect 13780 20896 13921 20924
rect 13780 20884 13786 20896
rect 13909 20893 13921 20896
rect 13955 20924 13967 20927
rect 14568 20924 14596 20964
rect 15105 20961 15117 20964
rect 15151 20961 15163 20995
rect 15105 20955 15163 20961
rect 13955 20896 14596 20924
rect 13955 20893 13967 20896
rect 13909 20887 13967 20893
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15212 20933 15240 21032
rect 17236 21032 20085 21060
rect 17236 21001 17264 21032
rect 20073 21029 20085 21032
rect 20119 21029 20131 21063
rect 20073 21023 20131 21029
rect 17221 20995 17279 21001
rect 17221 20961 17233 20995
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 17402 20952 17408 21004
rect 17460 20992 17466 21004
rect 18233 20995 18291 21001
rect 18233 20992 18245 20995
rect 17460 20964 18245 20992
rect 17460 20952 17466 20964
rect 18233 20961 18245 20964
rect 18279 20961 18291 20995
rect 18233 20955 18291 20961
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 20180 20992 20208 21100
rect 20349 21097 20361 21100
rect 20395 21097 20407 21131
rect 20349 21091 20407 21097
rect 20714 21088 20720 21140
rect 20772 21088 20778 21140
rect 21174 21128 21180 21140
rect 21008 21100 21180 21128
rect 20622 21060 20628 21072
rect 20456 21032 20628 21060
rect 20456 21001 20484 21032
rect 20622 21020 20628 21032
rect 20680 21020 20686 21072
rect 21008 21060 21036 21100
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 21821 21131 21879 21137
rect 21821 21097 21833 21131
rect 21867 21128 21879 21131
rect 22278 21128 22284 21140
rect 21867 21100 22284 21128
rect 21867 21097 21879 21100
rect 21821 21091 21879 21097
rect 22278 21088 22284 21100
rect 22336 21088 22342 21140
rect 23385 21131 23443 21137
rect 23385 21097 23397 21131
rect 23431 21128 23443 21131
rect 23934 21128 23940 21140
rect 23431 21100 23940 21128
rect 23431 21097 23443 21100
rect 23385 21091 23443 21097
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 24026 21088 24032 21140
rect 24084 21128 24090 21140
rect 24213 21131 24271 21137
rect 24213 21128 24225 21131
rect 24084 21100 24225 21128
rect 24084 21088 24090 21100
rect 24213 21097 24225 21100
rect 24259 21097 24271 21131
rect 24213 21091 24271 21097
rect 20732 21032 21036 21060
rect 19116 20964 20208 20992
rect 20441 20995 20499 21001
rect 19116 20952 19122 20964
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 17037 20927 17095 20933
rect 17037 20893 17049 20927
rect 17083 20924 17095 20927
rect 17310 20924 17316 20936
rect 17083 20896 17316 20924
rect 17083 20893 17095 20896
rect 17037 20887 17095 20893
rect 17310 20884 17316 20896
rect 17368 20884 17374 20936
rect 17494 20884 17500 20936
rect 17552 20924 17558 20936
rect 19444 20933 19472 20964
rect 20441 20961 20453 20995
rect 20487 20961 20499 20995
rect 20441 20955 20499 20961
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 17552 20896 18061 20924
rect 17552 20884 17558 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 14553 20859 14611 20865
rect 14553 20825 14565 20859
rect 14599 20856 14611 20859
rect 14599 20828 15240 20856
rect 14599 20825 14611 20828
rect 14553 20819 14611 20825
rect 15212 20800 15240 20828
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 19536 20856 19564 20887
rect 19702 20884 19708 20936
rect 19760 20884 19766 20936
rect 19886 20884 19892 20936
rect 19944 20884 19950 20936
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 19208 20828 19564 20856
rect 19996 20856 20024 20887
rect 20162 20884 20168 20936
rect 20220 20884 20226 20936
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20622 20884 20628 20936
rect 20680 20924 20686 20936
rect 20732 20924 20760 21032
rect 21008 20992 21036 21032
rect 21358 21020 21364 21072
rect 21416 21060 21422 21072
rect 21634 21060 21640 21072
rect 21416 21032 21640 21060
rect 21416 21020 21422 21032
rect 21634 21020 21640 21032
rect 21692 21020 21698 21072
rect 21177 20995 21235 21001
rect 21177 20992 21189 20995
rect 21008 20964 21189 20992
rect 21177 20961 21189 20964
rect 21223 20961 21235 20995
rect 21177 20955 21235 20961
rect 21545 20995 21603 21001
rect 21545 20961 21557 20995
rect 21591 20992 21603 20995
rect 23569 20995 23627 21001
rect 23569 20992 23581 20995
rect 21591 20964 23581 20992
rect 21591 20961 21603 20964
rect 21545 20955 21603 20961
rect 23569 20961 23581 20964
rect 23615 20961 23627 20995
rect 23569 20955 23627 20961
rect 23750 20952 23756 21004
rect 23808 20992 23814 21004
rect 24397 20995 24455 21001
rect 24397 20992 24409 20995
rect 23808 20964 24409 20992
rect 23808 20952 23814 20964
rect 24397 20961 24409 20964
rect 24443 20961 24455 20995
rect 24397 20955 24455 20961
rect 20680 20896 20760 20924
rect 20680 20884 20686 20896
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20926 21143 20927
rect 21266 20926 21272 20936
rect 21131 20898 21272 20926
rect 21131 20893 21143 20898
rect 21085 20887 21143 20893
rect 21266 20884 21272 20898
rect 21324 20884 21330 20936
rect 21358 20884 21364 20936
rect 21416 20884 21422 20936
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20924 21695 20927
rect 21726 20924 21732 20936
rect 21683 20896 21732 20924
rect 21683 20893 21695 20896
rect 21637 20887 21695 20893
rect 21726 20884 21732 20896
rect 21784 20884 21790 20936
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20924 21879 20927
rect 22465 20927 22523 20933
rect 21867 20896 22324 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 22296 20868 22324 20896
rect 22465 20893 22477 20927
rect 22511 20924 22523 20927
rect 22833 20927 22891 20933
rect 22833 20924 22845 20927
rect 22511 20896 22845 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 22833 20893 22845 20896
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 22922 20884 22928 20936
rect 22980 20924 22986 20936
rect 23017 20927 23075 20933
rect 23017 20924 23029 20927
rect 22980 20896 23029 20924
rect 22980 20884 22986 20896
rect 23017 20893 23029 20896
rect 23063 20893 23075 20927
rect 23017 20887 23075 20893
rect 23198 20884 23204 20936
rect 23256 20884 23262 20936
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 25222 20924 25228 20936
rect 23891 20896 25228 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 20714 20856 20720 20868
rect 19996 20828 20720 20856
rect 19208 20816 19214 20828
rect 20714 20816 20720 20828
rect 20772 20816 20778 20868
rect 21542 20856 21548 20868
rect 21473 20828 21548 20856
rect 12176 20760 13216 20788
rect 15194 20748 15200 20800
rect 15252 20748 15258 20800
rect 16666 20748 16672 20800
rect 16724 20748 16730 20800
rect 17129 20791 17187 20797
rect 17129 20757 17141 20791
rect 17175 20788 17187 20791
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 17175 20760 17509 20788
rect 17175 20757 17187 20760
rect 17129 20751 17187 20757
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 17497 20751 17555 20757
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18748 20760 18889 20788
rect 18748 20748 18754 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 18877 20751 18935 20757
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19521 20791 19579 20797
rect 19521 20788 19533 20791
rect 19484 20760 19533 20788
rect 19484 20748 19490 20760
rect 19521 20757 19533 20760
rect 19567 20757 19579 20791
rect 19521 20751 19579 20757
rect 19794 20748 19800 20800
rect 19852 20788 19858 20800
rect 21473 20788 21501 20828
rect 21542 20816 21548 20828
rect 21600 20856 21606 20868
rect 22097 20859 22155 20865
rect 22097 20856 22109 20859
rect 21600 20828 22109 20856
rect 21600 20816 21606 20828
rect 22097 20825 22109 20828
rect 22143 20825 22155 20859
rect 22097 20819 22155 20825
rect 22278 20816 22284 20868
rect 22336 20856 22342 20868
rect 22554 20856 22560 20868
rect 22336 20828 22560 20856
rect 22336 20816 22342 20828
rect 22554 20816 22560 20828
rect 22612 20816 22618 20868
rect 24670 20865 24676 20868
rect 23109 20859 23167 20865
rect 23109 20825 23121 20859
rect 23155 20825 23167 20859
rect 23109 20819 23167 20825
rect 24664 20819 24676 20865
rect 19852 20760 21501 20788
rect 19852 20748 19858 20760
rect 22002 20748 22008 20800
rect 22060 20748 22066 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23124 20788 23152 20819
rect 24670 20816 24676 20819
rect 24728 20816 24734 20868
rect 22704 20760 23152 20788
rect 22704 20748 22710 20760
rect 23658 20748 23664 20800
rect 23716 20788 23722 20800
rect 23753 20791 23811 20797
rect 23753 20788 23765 20791
rect 23716 20760 23765 20788
rect 23716 20748 23722 20760
rect 23753 20757 23765 20760
rect 23799 20757 23811 20791
rect 23753 20751 23811 20757
rect 25774 20748 25780 20800
rect 25832 20748 25838 20800
rect 1104 20698 26220 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 26220 20698
rect 1104 20624 26220 20646
rect 2041 20587 2099 20593
rect 2041 20553 2053 20587
rect 2087 20584 2099 20587
rect 2130 20584 2136 20596
rect 2087 20556 2136 20584
rect 2087 20553 2099 20556
rect 2041 20547 2099 20553
rect 2130 20544 2136 20556
rect 2188 20544 2194 20596
rect 2314 20544 2320 20596
rect 2372 20544 2378 20596
rect 2406 20544 2412 20596
rect 2464 20584 2470 20596
rect 2464 20556 5396 20584
rect 2464 20544 2470 20556
rect 2774 20476 2780 20528
rect 2832 20516 2838 20528
rect 2929 20519 2987 20525
rect 2929 20516 2941 20519
rect 2832 20488 2941 20516
rect 2832 20476 2838 20488
rect 2929 20485 2941 20488
rect 2975 20485 2987 20519
rect 2929 20479 2987 20485
rect 3145 20519 3203 20525
rect 3145 20485 3157 20519
rect 3191 20516 3203 20519
rect 3234 20516 3240 20528
rect 3191 20488 3240 20516
rect 3191 20485 3203 20488
rect 3145 20479 3203 20485
rect 3234 20476 3240 20488
rect 3292 20516 3298 20528
rect 3421 20519 3479 20525
rect 3421 20516 3433 20519
rect 3292 20488 3433 20516
rect 3292 20476 3298 20488
rect 3421 20485 3433 20488
rect 3467 20485 3479 20519
rect 3421 20479 3479 20485
rect 3786 20476 3792 20528
rect 3844 20476 3850 20528
rect 4062 20476 4068 20528
rect 4120 20516 4126 20528
rect 5368 20525 5396 20556
rect 7374 20544 7380 20596
rect 7432 20584 7438 20596
rect 9306 20584 9312 20596
rect 7432 20556 9312 20584
rect 7432 20544 7438 20556
rect 9306 20544 9312 20556
rect 9364 20584 9370 20596
rect 9364 20556 9812 20584
rect 9364 20544 9370 20556
rect 5353 20519 5411 20525
rect 4120 20488 4844 20516
rect 4120 20476 4126 20488
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 1780 20312 1808 20411
rect 1946 20408 1952 20460
rect 2004 20408 2010 20460
rect 2409 20451 2467 20457
rect 2409 20417 2421 20451
rect 2455 20448 2467 20451
rect 2498 20448 2504 20460
rect 2455 20420 2504 20448
rect 2455 20417 2467 20420
rect 2409 20411 2467 20417
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 2682 20408 2688 20460
rect 2740 20408 2746 20460
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 2200 20383 2258 20389
rect 2200 20380 2212 20383
rect 1903 20352 2212 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 2200 20349 2212 20352
rect 2246 20349 2258 20383
rect 2200 20343 2258 20349
rect 3237 20383 3295 20389
rect 3237 20349 3249 20383
rect 3283 20380 3295 20383
rect 3418 20380 3424 20392
rect 3283 20352 3424 20380
rect 3283 20349 3295 20352
rect 3237 20343 3295 20349
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 2777 20315 2835 20321
rect 2777 20312 2789 20315
rect 1780 20284 2789 20312
rect 2777 20281 2789 20284
rect 2823 20312 2835 20315
rect 2866 20312 2872 20324
rect 2823 20284 2872 20312
rect 2823 20281 2835 20284
rect 2777 20275 2835 20281
rect 2866 20272 2872 20284
rect 2924 20272 2930 20324
rect 2222 20204 2228 20256
rect 2280 20244 2286 20256
rect 2961 20247 3019 20253
rect 2961 20244 2973 20247
rect 2280 20216 2973 20244
rect 2280 20204 2286 20216
rect 2961 20213 2973 20216
rect 3007 20244 3019 20247
rect 3528 20244 3556 20411
rect 3602 20408 3608 20460
rect 3660 20408 3666 20460
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4522 20448 4528 20460
rect 4479 20420 4528 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 4614 20408 4620 20460
rect 4672 20408 4678 20460
rect 4706 20408 4712 20460
rect 4764 20408 4770 20460
rect 4816 20457 4844 20488
rect 5353 20485 5365 20519
rect 5399 20516 5411 20519
rect 5399 20488 6408 20516
rect 5399 20485 5411 20488
rect 5353 20479 5411 20485
rect 6380 20457 6408 20488
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 8665 20519 8723 20525
rect 8665 20516 8677 20519
rect 8352 20488 8677 20516
rect 8352 20476 8358 20488
rect 8665 20485 8677 20488
rect 8711 20516 8723 20519
rect 9030 20516 9036 20528
rect 8711 20488 9036 20516
rect 8711 20485 8723 20488
rect 8665 20479 8723 20485
rect 9030 20476 9036 20488
rect 9088 20476 9094 20528
rect 9122 20476 9128 20528
rect 9180 20516 9186 20528
rect 9180 20488 9628 20516
rect 9180 20476 9186 20488
rect 9600 20457 9628 20488
rect 9784 20457 9812 20556
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12584 20556 12848 20584
rect 12584 20544 12590 20556
rect 12434 20476 12440 20528
rect 12492 20516 12498 20528
rect 12492 20488 12572 20516
rect 12492 20476 12498 20488
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 6181 20451 6239 20457
rect 6181 20417 6193 20451
rect 6227 20417 6239 20451
rect 6181 20411 6239 20417
rect 6365 20451 6423 20457
rect 6365 20417 6377 20451
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 9493 20451 9551 20457
rect 9493 20417 9505 20451
rect 9539 20417 9551 20451
rect 9493 20411 9551 20417
rect 9585 20451 9643 20457
rect 9585 20417 9597 20451
rect 9631 20417 9643 20451
rect 9585 20411 9643 20417
rect 9769 20451 9827 20457
rect 9769 20417 9781 20451
rect 9815 20417 9827 20451
rect 12544 20448 12572 20488
rect 12618 20476 12624 20528
rect 12676 20525 12682 20528
rect 12676 20516 12688 20525
rect 12820 20516 12848 20556
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12952 20556 13001 20584
rect 12952 20544 12958 20556
rect 12989 20553 13001 20556
rect 13035 20553 13047 20587
rect 12989 20547 13047 20553
rect 13357 20587 13415 20593
rect 13357 20553 13369 20587
rect 13403 20584 13415 20587
rect 13814 20584 13820 20596
rect 13403 20556 13820 20584
rect 13403 20553 13415 20556
rect 13357 20547 13415 20553
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 13998 20544 14004 20596
rect 14056 20544 14062 20596
rect 15194 20544 15200 20596
rect 15252 20544 15258 20596
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20584 15715 20587
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 15703 20556 16681 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 16669 20553 16681 20556
rect 16715 20584 16727 20587
rect 17402 20584 17408 20596
rect 16715 20556 17408 20584
rect 16715 20553 16727 20556
rect 16669 20547 16727 20553
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 18141 20587 18199 20593
rect 18141 20553 18153 20587
rect 18187 20553 18199 20587
rect 19794 20584 19800 20596
rect 18141 20547 18199 20553
rect 18340 20556 19800 20584
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 12676 20488 12721 20516
rect 12820 20488 13737 20516
rect 12676 20479 12688 20488
rect 13725 20485 13737 20488
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 13909 20519 13967 20525
rect 13909 20485 13921 20519
rect 13955 20516 13967 20519
rect 14090 20516 14096 20528
rect 13955 20488 14096 20516
rect 13955 20485 13967 20488
rect 13909 20479 13967 20485
rect 12676 20476 12682 20479
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 15010 20516 15016 20528
rect 14200 20488 15016 20516
rect 12544 20420 13032 20448
rect 9769 20411 9827 20417
rect 4540 20380 4568 20408
rect 5074 20380 5080 20392
rect 4540 20352 5080 20380
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 6196 20380 6224 20411
rect 9508 20380 9536 20411
rect 10502 20380 10508 20392
rect 6196 20352 10508 20380
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 12894 20340 12900 20392
rect 12952 20340 12958 20392
rect 13004 20380 13032 20420
rect 13170 20408 13176 20460
rect 13228 20408 13234 20460
rect 13446 20408 13452 20460
rect 13504 20408 13510 20460
rect 13538 20408 13544 20460
rect 13596 20448 13602 20460
rect 14200 20457 14228 20488
rect 15010 20476 15016 20488
rect 15068 20476 15074 20528
rect 17804 20519 17862 20525
rect 17804 20485 17816 20519
rect 17850 20516 17862 20519
rect 18156 20516 18184 20547
rect 17850 20488 18184 20516
rect 17850 20485 17862 20488
rect 17804 20479 17862 20485
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13596 20420 14197 20448
rect 13596 20408 13602 20420
rect 14185 20417 14197 20420
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 14366 20408 14372 20460
rect 14424 20408 14430 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 15565 20451 15623 20457
rect 15565 20448 15577 20451
rect 15436 20420 15577 20448
rect 15436 20408 15442 20420
rect 15565 20417 15577 20420
rect 15611 20417 15623 20451
rect 17310 20448 17316 20460
rect 15565 20411 15623 20417
rect 15856 20420 17316 20448
rect 14384 20380 14412 20408
rect 13004 20352 14412 20380
rect 14458 20340 14464 20392
rect 14516 20340 14522 20392
rect 15856 20389 15884 20420
rect 17310 20408 17316 20420
rect 17368 20408 17374 20460
rect 18340 20457 18368 20556
rect 19794 20544 19800 20556
rect 19852 20544 19858 20596
rect 20622 20544 20628 20596
rect 20680 20584 20686 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20680 20556 21005 20584
rect 20680 20544 20686 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 21358 20544 21364 20596
rect 21416 20544 21422 20596
rect 22922 20584 22928 20596
rect 22848 20556 22928 20584
rect 18509 20519 18567 20525
rect 18509 20485 18521 20519
rect 18555 20516 18567 20519
rect 18785 20519 18843 20525
rect 18785 20516 18797 20519
rect 18555 20488 18797 20516
rect 18555 20485 18567 20488
rect 18509 20479 18567 20485
rect 18785 20485 18797 20488
rect 18831 20485 18843 20519
rect 19426 20516 19432 20528
rect 18785 20479 18843 20485
rect 18892 20488 19432 20516
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20417 18475 20451
rect 18417 20411 18475 20417
rect 15841 20383 15899 20389
rect 15841 20349 15853 20383
rect 15887 20349 15899 20383
rect 15841 20343 15899 20349
rect 18046 20340 18052 20392
rect 18104 20340 18110 20392
rect 18432 20380 18460 20411
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 18892 20380 18920 20488
rect 19426 20476 19432 20488
rect 19484 20476 19490 20528
rect 22186 20516 22192 20528
rect 21376 20488 22192 20516
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 18432 20352 18920 20380
rect 13354 20312 13360 20324
rect 12912 20284 13360 20312
rect 3007 20216 3556 20244
rect 5077 20247 5135 20253
rect 3007 20213 3019 20216
rect 2961 20207 3019 20213
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5166 20244 5172 20256
rect 5123 20216 5172 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 9585 20247 9643 20253
rect 9585 20244 9597 20247
rect 8720 20216 9597 20244
rect 8720 20204 8726 20216
rect 9585 20213 9597 20216
rect 9631 20213 9643 20247
rect 9585 20207 9643 20213
rect 11517 20247 11575 20253
rect 11517 20213 11529 20247
rect 11563 20244 11575 20247
rect 12526 20244 12532 20256
rect 11563 20216 12532 20244
rect 11563 20213 11575 20216
rect 11517 20207 11575 20213
rect 12526 20204 12532 20216
rect 12584 20244 12590 20256
rect 12912 20244 12940 20284
rect 13354 20272 13360 20284
rect 13412 20272 13418 20324
rect 15105 20315 15163 20321
rect 15105 20281 15117 20315
rect 15151 20312 15163 20315
rect 15286 20312 15292 20324
rect 15151 20284 15292 20312
rect 15151 20281 15163 20284
rect 15105 20275 15163 20281
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 18984 20312 19012 20411
rect 19076 20380 19104 20411
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19702 20448 19708 20460
rect 19392 20420 19708 20448
rect 19392 20408 19398 20420
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 20533 20451 20591 20457
rect 20533 20448 20545 20451
rect 20220 20420 20545 20448
rect 20220 20408 20226 20420
rect 20533 20417 20545 20420
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21177 20451 21235 20457
rect 20947 20420 21036 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 19886 20380 19892 20392
rect 19076 20352 19892 20380
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 19794 20312 19800 20324
rect 18984 20284 19800 20312
rect 19794 20272 19800 20284
rect 19852 20272 19858 20324
rect 20530 20272 20536 20324
rect 20588 20312 20594 20324
rect 20640 20312 20668 20411
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 20809 20383 20867 20389
rect 20809 20380 20821 20383
rect 20772 20352 20821 20380
rect 20772 20340 20778 20352
rect 20809 20349 20821 20352
rect 20855 20349 20867 20383
rect 20809 20343 20867 20349
rect 20588 20284 20668 20312
rect 21008 20312 21036 20420
rect 21177 20417 21189 20451
rect 21223 20446 21235 20451
rect 21376 20448 21404 20488
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 22848 20525 22876 20556
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 23106 20544 23112 20596
rect 23164 20584 23170 20596
rect 23164 20556 23612 20584
rect 23164 20544 23170 20556
rect 22833 20519 22891 20525
rect 22833 20485 22845 20519
rect 22879 20516 22891 20519
rect 23477 20519 23535 20525
rect 23477 20516 23489 20519
rect 22879 20488 23489 20516
rect 22879 20485 22891 20488
rect 22833 20479 22891 20485
rect 23477 20485 23489 20488
rect 23523 20485 23535 20519
rect 23584 20516 23612 20556
rect 23658 20544 23664 20596
rect 23716 20584 23722 20596
rect 23845 20587 23903 20593
rect 23845 20584 23857 20587
rect 23716 20556 23857 20584
rect 23716 20544 23722 20556
rect 23845 20553 23857 20556
rect 23891 20553 23903 20587
rect 23845 20547 23903 20553
rect 24670 20544 24676 20596
rect 24728 20544 24734 20596
rect 24949 20587 25007 20593
rect 24949 20553 24961 20587
rect 24995 20584 25007 20587
rect 25590 20584 25596 20596
rect 24995 20556 25596 20584
rect 24995 20553 25007 20556
rect 24949 20547 25007 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 24305 20519 24363 20525
rect 23584 20488 23704 20516
rect 23477 20479 23535 20485
rect 21284 20446 21404 20448
rect 21223 20420 21404 20446
rect 21453 20451 21511 20457
rect 21223 20418 21312 20420
rect 21223 20417 21235 20418
rect 21177 20411 21235 20417
rect 21453 20417 21465 20451
rect 21499 20448 21511 20451
rect 21634 20448 21640 20460
rect 21499 20420 21640 20448
rect 21499 20417 21511 20420
rect 21453 20411 21511 20417
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 21910 20448 21916 20460
rect 21867 20420 21916 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 21910 20408 21916 20420
rect 21968 20408 21974 20460
rect 22005 20451 22063 20457
rect 22005 20417 22017 20451
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 21082 20340 21088 20392
rect 21140 20380 21146 20392
rect 22020 20380 22048 20411
rect 22094 20408 22100 20460
rect 22152 20408 22158 20460
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 21140 20352 22048 20380
rect 21140 20340 21146 20352
rect 22186 20340 22192 20392
rect 22244 20340 22250 20392
rect 21266 20312 21272 20324
rect 21008 20284 21272 20312
rect 20588 20272 20594 20284
rect 12584 20216 12940 20244
rect 12584 20204 12590 20216
rect 12986 20204 12992 20256
rect 13044 20244 13050 20256
rect 13446 20244 13452 20256
rect 13044 20216 13452 20244
rect 13044 20204 13050 20216
rect 13446 20204 13452 20216
rect 13504 20244 13510 20256
rect 13541 20247 13599 20253
rect 13541 20244 13553 20247
rect 13504 20216 13553 20244
rect 13504 20204 13510 20216
rect 13541 20213 13553 20216
rect 13587 20213 13599 20247
rect 13541 20207 13599 20213
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 15194 20244 15200 20256
rect 14332 20216 15200 20244
rect 14332 20204 14338 20216
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 20346 20204 20352 20256
rect 20404 20204 20410 20256
rect 20640 20244 20668 20284
rect 21266 20272 21272 20284
rect 21324 20312 21330 20324
rect 22002 20312 22008 20324
rect 21324 20284 22008 20312
rect 21324 20272 21330 20284
rect 22002 20272 22008 20284
rect 22060 20312 22066 20324
rect 22388 20312 22416 20411
rect 22462 20408 22468 20460
rect 22520 20448 22526 20460
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22520 20420 22661 20448
rect 22520 20408 22526 20420
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22649 20411 22707 20417
rect 22848 20420 22937 20448
rect 22848 20392 22876 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23106 20448 23112 20460
rect 23063 20420 23112 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23290 20408 23296 20460
rect 23348 20408 23354 20460
rect 23566 20408 23572 20460
rect 23624 20408 23630 20460
rect 23676 20457 23704 20488
rect 24305 20485 24317 20519
rect 24351 20516 24363 20519
rect 25041 20519 25099 20525
rect 25041 20516 25053 20519
rect 24351 20488 25053 20516
rect 24351 20485 24363 20488
rect 24305 20479 24363 20485
rect 25041 20485 25053 20488
rect 25087 20485 25099 20519
rect 25041 20479 25099 20485
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 25685 20451 25743 20457
rect 25685 20448 25697 20451
rect 24811 20420 25697 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 25685 20417 25697 20420
rect 25731 20448 25743 20451
rect 25774 20448 25780 20460
rect 25731 20420 25780 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 22830 20340 22836 20392
rect 22888 20340 22894 20392
rect 24029 20383 24087 20389
rect 24029 20380 24041 20383
rect 23124 20352 24041 20380
rect 22060 20284 22416 20312
rect 22557 20315 22615 20321
rect 22060 20272 22066 20284
rect 22557 20281 22569 20315
rect 22603 20312 22615 20315
rect 23124 20312 23152 20352
rect 24029 20349 24041 20352
rect 24075 20349 24087 20383
rect 24029 20343 24087 20349
rect 24213 20383 24271 20389
rect 24213 20349 24225 20383
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 22603 20284 23152 20312
rect 23201 20315 23259 20321
rect 22603 20281 22615 20284
rect 22557 20275 22615 20281
rect 23201 20281 23213 20315
rect 23247 20312 23259 20315
rect 24228 20312 24256 20343
rect 23247 20284 24256 20312
rect 23247 20281 23259 20284
rect 23201 20275 23259 20281
rect 23106 20244 23112 20256
rect 20640 20216 23112 20244
rect 23106 20204 23112 20216
rect 23164 20204 23170 20256
rect 1104 20154 26220 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 26220 20154
rect 1104 20080 26220 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2004 20012 2973 20040
rect 2004 20000 2010 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 2961 20003 3019 20009
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 3786 20040 3792 20052
rect 3292 20012 3792 20040
rect 3292 20000 3298 20012
rect 3786 20000 3792 20012
rect 3844 20040 3850 20052
rect 4249 20043 4307 20049
rect 4249 20040 4261 20043
rect 3844 20012 4261 20040
rect 3844 20000 3850 20012
rect 4249 20009 4261 20012
rect 4295 20009 4307 20043
rect 4249 20003 4307 20009
rect 6365 20043 6423 20049
rect 6365 20009 6377 20043
rect 6411 20040 6423 20043
rect 6822 20040 6828 20052
rect 6411 20012 6828 20040
rect 6411 20009 6423 20012
rect 6365 20003 6423 20009
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 8386 20000 8392 20052
rect 8444 20000 8450 20052
rect 14185 20043 14243 20049
rect 14185 20009 14197 20043
rect 14231 20040 14243 20043
rect 14458 20040 14464 20052
rect 14231 20012 14464 20040
rect 14231 20009 14243 20012
rect 14185 20003 14243 20009
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 17037 20043 17095 20049
rect 17037 20009 17049 20043
rect 17083 20040 17095 20043
rect 17126 20040 17132 20052
rect 17083 20012 17132 20040
rect 17083 20009 17095 20012
rect 17037 20003 17095 20009
rect 17126 20000 17132 20012
rect 17184 20040 17190 20052
rect 17494 20040 17500 20052
rect 17184 20012 17500 20040
rect 17184 20000 17190 20012
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19484 20012 20760 20040
rect 19484 20000 19490 20012
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19941 4675 19975
rect 8294 19972 8300 19984
rect 4617 19935 4675 19941
rect 8128 19944 8300 19972
rect 3602 19904 3608 19916
rect 2792 19876 3608 19904
rect 2792 19848 2820 19876
rect 3602 19864 3608 19876
rect 3660 19864 3666 19916
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4341 19907 4399 19913
rect 4341 19904 4353 19907
rect 4120 19876 4353 19904
rect 4120 19864 4126 19876
rect 4341 19873 4353 19876
rect 4387 19873 4399 19907
rect 4632 19904 4660 19935
rect 4632 19876 5396 19904
rect 4341 19867 4399 19873
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 2774 19836 2780 19848
rect 2731 19808 2780 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19836 3019 19839
rect 3234 19836 3240 19848
rect 3007 19808 3240 19836
rect 3007 19805 3019 19808
rect 2961 19799 3019 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 3936 19808 4261 19836
rect 3936 19796 3942 19808
rect 4249 19805 4261 19808
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4672 19808 4905 19836
rect 4672 19796 4678 19808
rect 4893 19805 4905 19808
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 5074 19796 5080 19848
rect 5132 19796 5138 19848
rect 5166 19796 5172 19848
rect 5224 19796 5230 19848
rect 5368 19845 5396 19876
rect 5644 19876 6500 19904
rect 5644 19848 5672 19876
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19836 5595 19839
rect 5626 19836 5632 19848
rect 5583 19808 5632 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 5460 19768 5488 19799
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 6472 19845 6500 19876
rect 7742 19864 7748 19916
rect 7800 19864 7806 19916
rect 8128 19913 8156 19944
rect 8294 19932 8300 19944
rect 8352 19972 8358 19984
rect 8478 19972 8484 19984
rect 8352 19944 8484 19972
rect 8352 19932 8358 19944
rect 8478 19932 8484 19944
rect 8536 19932 8542 19984
rect 19334 19932 19340 19984
rect 19392 19972 19398 19984
rect 20257 19975 20315 19981
rect 20257 19972 20269 19975
rect 19392 19944 20269 19972
rect 19392 19932 19398 19944
rect 20257 19941 20269 19944
rect 20303 19941 20315 19975
rect 20257 19935 20315 19941
rect 8113 19907 8171 19913
rect 8113 19873 8125 19907
rect 8159 19873 8171 19907
rect 8938 19904 8944 19916
rect 8113 19867 8171 19873
rect 8496 19876 8944 19904
rect 8496 19848 8524 19876
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 15654 19904 15660 19916
rect 15611 19876 15660 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 19058 19864 19064 19916
rect 19116 19904 19122 19916
rect 20349 19907 20407 19913
rect 20349 19904 20361 19907
rect 19116 19876 20361 19904
rect 19116 19864 19122 19876
rect 20349 19873 20361 19876
rect 20395 19873 20407 19907
rect 20349 19867 20407 19873
rect 20625 19907 20683 19913
rect 20625 19873 20637 19907
rect 20671 19873 20683 19907
rect 20625 19867 20683 19873
rect 6089 19839 6147 19845
rect 6089 19836 6101 19839
rect 5776 19808 6101 19836
rect 5776 19796 5782 19808
rect 6089 19805 6101 19808
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 6457 19839 6515 19845
rect 6457 19805 6469 19839
rect 6503 19836 6515 19839
rect 6733 19839 6791 19845
rect 6733 19836 6745 19839
rect 6503 19808 6745 19836
rect 6503 19805 6515 19808
rect 6457 19799 6515 19805
rect 6733 19805 6745 19808
rect 6779 19805 6791 19839
rect 6733 19799 6791 19805
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8662 19796 8668 19848
rect 8720 19796 8726 19848
rect 9030 19796 9036 19848
rect 9088 19796 9094 19848
rect 10502 19796 10508 19848
rect 10560 19836 10566 19848
rect 11054 19836 11060 19848
rect 10560 19808 11060 19836
rect 10560 19796 10566 19808
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 11333 19839 11391 19845
rect 11333 19805 11345 19839
rect 11379 19836 11391 19839
rect 11514 19836 11520 19848
rect 11379 19808 11520 19836
rect 11379 19805 11391 19808
rect 11333 19799 11391 19805
rect 11514 19796 11520 19808
rect 11572 19836 11578 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11572 19808 11713 19836
rect 11572 19796 11578 19808
rect 11701 19805 11713 19808
rect 11747 19836 11759 19839
rect 12066 19836 12072 19848
rect 11747 19808 12072 19836
rect 11747 19805 11759 19808
rect 11701 19799 11759 19805
rect 12066 19796 12072 19808
rect 12124 19836 12130 19848
rect 12894 19836 12900 19848
rect 12124 19808 12900 19836
rect 12124 19796 12130 19808
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 14090 19836 14096 19848
rect 13955 19808 14096 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 6549 19771 6607 19777
rect 6549 19768 6561 19771
rect 5460 19740 6561 19768
rect 6549 19737 6561 19740
rect 6595 19768 6607 19771
rect 6822 19768 6828 19780
rect 6595 19740 6828 19768
rect 6595 19737 6607 19740
rect 6549 19731 6607 19737
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 8230 19771 8288 19777
rect 8230 19737 8242 19771
rect 8276 19768 8288 19771
rect 8573 19771 8631 19777
rect 8573 19768 8585 19771
rect 8276 19740 8585 19768
rect 8276 19737 8288 19740
rect 8230 19731 8288 19737
rect 8573 19737 8585 19740
rect 8619 19737 8631 19771
rect 8573 19731 8631 19737
rect 11422 19728 11428 19780
rect 11480 19768 11486 19780
rect 11882 19768 11888 19780
rect 11480 19740 11888 19768
rect 11480 19728 11486 19740
rect 11882 19728 11888 19740
rect 11940 19768 11946 19780
rect 13740 19768 13768 19799
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 15924 19839 15982 19845
rect 15924 19805 15936 19839
rect 15970 19836 15982 19839
rect 16666 19836 16672 19848
rect 15970 19808 16672 19836
rect 15970 19805 15982 19808
rect 15924 19799 15982 19805
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 18046 19796 18052 19848
rect 18104 19836 18110 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18104 19808 18889 19836
rect 18104 19796 18110 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 19242 19796 19248 19848
rect 19300 19796 19306 19848
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 19944 19808 20177 19836
rect 19944 19796 19950 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19836 20499 19839
rect 20640 19836 20668 19867
rect 20487 19808 20668 19836
rect 20732 19836 20760 20012
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 21910 20040 21916 20052
rect 20864 20012 21916 20040
rect 20864 20000 20870 20012
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 22186 20000 22192 20052
rect 22244 20000 22250 20052
rect 20990 19972 20996 19984
rect 20824 19944 20996 19972
rect 20824 19913 20852 19944
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 21358 19932 21364 19984
rect 21416 19972 21422 19984
rect 22097 19975 22155 19981
rect 21416 19944 21772 19972
rect 21416 19932 21422 19944
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19873 20867 19907
rect 20809 19867 20867 19873
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19904 20959 19907
rect 21174 19904 21180 19916
rect 20947 19876 21180 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 20990 19836 20996 19848
rect 20732 19808 20996 19836
rect 20487 19805 20499 19808
rect 20441 19799 20499 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19836 21143 19839
rect 21131 19808 21220 19836
rect 21131 19805 21143 19808
rect 21085 19799 21143 19805
rect 11940 19740 13768 19768
rect 11940 19728 11946 19740
rect 14826 19728 14832 19780
rect 14884 19768 14890 19780
rect 15298 19771 15356 19777
rect 15298 19768 15310 19771
rect 14884 19740 15310 19768
rect 14884 19728 14890 19740
rect 15298 19737 15310 19740
rect 15344 19737 15356 19771
rect 15298 19731 15356 19737
rect 18632 19771 18690 19777
rect 18632 19737 18644 19771
rect 18678 19768 18690 19771
rect 19981 19771 20039 19777
rect 19981 19768 19993 19771
rect 18678 19740 19993 19768
rect 18678 19737 18690 19740
rect 18632 19731 18690 19737
rect 19981 19737 19993 19740
rect 20027 19737 20039 19771
rect 19981 19731 20039 19737
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 2777 19703 2835 19709
rect 2777 19700 2789 19703
rect 2280 19672 2789 19700
rect 2280 19660 2286 19672
rect 2777 19669 2789 19672
rect 2823 19669 2835 19703
rect 2777 19663 2835 19669
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5626 19700 5632 19712
rect 5123 19672 5632 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 5810 19660 5816 19712
rect 5868 19660 5874 19712
rect 5902 19660 5908 19712
rect 5960 19660 5966 19712
rect 6914 19660 6920 19712
rect 6972 19660 6978 19712
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8662 19700 8668 19712
rect 8067 19672 8668 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 13814 19660 13820 19712
rect 13872 19660 13878 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 18322 19700 18328 19712
rect 17543 19672 18328 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18322 19660 18328 19672
rect 18380 19700 18386 19712
rect 19242 19700 19248 19712
rect 18380 19672 19248 19700
rect 18380 19660 18386 19672
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19889 19703 19947 19709
rect 19889 19669 19901 19703
rect 19935 19700 19947 19703
rect 21192 19700 21220 19808
rect 21358 19796 21364 19848
rect 21416 19836 21422 19848
rect 21634 19836 21640 19848
rect 21416 19808 21640 19836
rect 21416 19796 21422 19808
rect 21634 19796 21640 19808
rect 21692 19796 21698 19848
rect 21744 19845 21772 19944
rect 22097 19941 22109 19975
rect 22143 19972 22155 19975
rect 23290 19972 23296 19984
rect 22143 19944 23296 19972
rect 22143 19941 22155 19944
rect 22097 19935 22155 19941
rect 23290 19932 23296 19944
rect 23348 19932 23354 19984
rect 22462 19864 22468 19916
rect 22520 19904 22526 19916
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 22520 19876 24961 19904
rect 22520 19864 22526 19876
rect 24949 19873 24961 19876
rect 24995 19873 25007 19907
rect 24949 19867 25007 19873
rect 21729 19839 21787 19845
rect 21729 19805 21741 19839
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19836 21971 19839
rect 22094 19836 22100 19848
rect 21959 19808 22100 19836
rect 21959 19805 21971 19808
rect 21913 19799 21971 19805
rect 22094 19796 22100 19808
rect 22152 19836 22158 19848
rect 22278 19836 22284 19848
rect 22152 19808 22284 19836
rect 22152 19796 22158 19808
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 22554 19796 22560 19848
rect 22612 19796 22618 19848
rect 23934 19796 23940 19848
rect 23992 19796 23998 19848
rect 25314 19796 25320 19848
rect 25372 19836 25378 19848
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25372 19808 25789 19836
rect 25372 19796 25378 19808
rect 25777 19805 25789 19808
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 22370 19728 22376 19780
rect 22428 19728 22434 19780
rect 24765 19771 24823 19777
rect 24765 19737 24777 19771
rect 24811 19768 24823 19771
rect 25225 19771 25283 19777
rect 25225 19768 25237 19771
rect 24811 19740 25237 19768
rect 24811 19737 24823 19740
rect 24765 19731 24823 19737
rect 25225 19737 25237 19740
rect 25271 19737 25283 19771
rect 25225 19731 25283 19737
rect 19935 19672 21220 19700
rect 19935 19669 19947 19672
rect 19889 19663 19947 19669
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21818 19700 21824 19712
rect 21324 19672 21824 19700
rect 21324 19660 21330 19672
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 23842 19700 23848 19712
rect 23624 19672 23848 19700
rect 23624 19660 23630 19672
rect 23842 19660 23848 19672
rect 23900 19660 23906 19712
rect 24118 19660 24124 19712
rect 24176 19660 24182 19712
rect 24394 19660 24400 19712
rect 24452 19660 24458 19712
rect 24486 19660 24492 19712
rect 24544 19700 24550 19712
rect 24857 19703 24915 19709
rect 24857 19700 24869 19703
rect 24544 19672 24869 19700
rect 24544 19660 24550 19672
rect 24857 19669 24869 19672
rect 24903 19669 24915 19703
rect 24857 19663 24915 19669
rect 1104 19610 26220 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 26220 19610
rect 1104 19536 26220 19558
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 12492 19468 12909 19496
rect 12492 19456 12498 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 13906 19456 13912 19508
rect 13964 19456 13970 19508
rect 14369 19499 14427 19505
rect 14369 19465 14381 19499
rect 14415 19496 14427 19499
rect 14458 19496 14464 19508
rect 14415 19468 14464 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14826 19456 14832 19508
rect 14884 19456 14890 19508
rect 19058 19456 19064 19508
rect 19116 19456 19122 19508
rect 20990 19456 20996 19508
rect 21048 19496 21054 19508
rect 21243 19499 21301 19505
rect 21243 19496 21255 19499
rect 21048 19468 21255 19496
rect 21048 19456 21054 19468
rect 21243 19465 21255 19468
rect 21289 19465 21301 19499
rect 22186 19496 22192 19508
rect 21243 19459 21301 19465
rect 21468 19468 22192 19496
rect 2314 19388 2320 19440
rect 2372 19428 2378 19440
rect 3142 19428 3148 19440
rect 2372 19400 2728 19428
rect 2372 19388 2378 19400
rect 2222 19320 2228 19372
rect 2280 19320 2286 19372
rect 2700 19369 2728 19400
rect 2792 19400 3148 19428
rect 2685 19363 2743 19369
rect 2685 19329 2697 19363
rect 2731 19360 2743 19363
rect 2792 19360 2820 19400
rect 3142 19388 3148 19400
rect 3200 19388 3206 19440
rect 3252 19400 5672 19428
rect 2731 19332 2820 19360
rect 2869 19363 2927 19369
rect 2731 19329 2743 19332
rect 2685 19323 2743 19329
rect 2869 19329 2881 19363
rect 2915 19360 2927 19363
rect 3252 19360 3280 19400
rect 2915 19332 3280 19360
rect 2915 19329 2927 19332
rect 2869 19323 2927 19329
rect 3786 19320 3792 19372
rect 3844 19320 3850 19372
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 4120 19332 4445 19360
rect 4120 19320 4126 19332
rect 4433 19329 4445 19332
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 4764 19332 5549 19360
rect 4764 19320 4770 19332
rect 5537 19329 5549 19332
rect 5583 19329 5595 19363
rect 5537 19323 5595 19329
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2774 19292 2780 19304
rect 2363 19264 2780 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 3878 19252 3884 19304
rect 3936 19252 3942 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4614 19292 4620 19304
rect 4571 19264 4620 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 4157 19227 4215 19233
rect 4157 19193 4169 19227
rect 4203 19224 4215 19227
rect 4724 19224 4752 19320
rect 4203 19196 4752 19224
rect 5644 19224 5672 19400
rect 5810 19388 5816 19440
rect 5868 19428 5874 19440
rect 5868 19400 6500 19428
rect 5868 19388 5874 19400
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19360 5779 19363
rect 5902 19360 5908 19372
rect 5767 19332 5908 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 6472 19369 6500 19400
rect 7834 19388 7840 19440
rect 7892 19428 7898 19440
rect 8202 19428 8208 19440
rect 7892 19400 8208 19428
rect 7892 19388 7898 19400
rect 8202 19388 8208 19400
rect 8260 19428 8266 19440
rect 9033 19431 9091 19437
rect 9033 19428 9045 19431
rect 8260 19400 9045 19428
rect 8260 19388 8266 19400
rect 9033 19397 9045 19400
rect 9079 19397 9091 19431
rect 9033 19391 9091 19397
rect 10965 19431 11023 19437
rect 10965 19397 10977 19431
rect 11011 19428 11023 19431
rect 11762 19431 11820 19437
rect 11762 19428 11774 19431
rect 11011 19400 11774 19428
rect 11011 19397 11023 19400
rect 10965 19391 11023 19397
rect 11762 19397 11774 19400
rect 11808 19397 11820 19431
rect 19426 19428 19432 19440
rect 11762 19391 11820 19397
rect 18892 19400 19432 19428
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6052 19332 6377 19360
rect 6052 19320 6058 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6458 19363 6516 19369
rect 6458 19329 6470 19363
rect 6504 19329 6516 19363
rect 6458 19323 6516 19329
rect 6546 19320 6552 19372
rect 6604 19360 6610 19372
rect 6914 19369 6920 19372
rect 6641 19363 6699 19369
rect 6641 19360 6653 19363
rect 6604 19332 6653 19360
rect 6604 19320 6610 19332
rect 6641 19329 6653 19332
rect 6687 19329 6699 19363
rect 6641 19323 6699 19329
rect 6733 19363 6791 19369
rect 6733 19329 6745 19363
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 6871 19363 6920 19369
rect 6871 19329 6883 19363
rect 6917 19329 6920 19363
rect 6871 19323 6920 19329
rect 5920 19292 5948 19320
rect 6748 19292 6776 19323
rect 6914 19320 6920 19323
rect 6972 19320 6978 19372
rect 8386 19320 8392 19372
rect 8444 19320 8450 19372
rect 10689 19363 10747 19369
rect 10689 19329 10701 19363
rect 10735 19360 10747 19363
rect 11422 19360 11428 19372
rect 10735 19332 11428 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 11422 19320 11428 19332
rect 11480 19320 11486 19372
rect 11514 19320 11520 19372
rect 11572 19320 11578 19372
rect 14090 19320 14096 19372
rect 14148 19360 14154 19372
rect 14461 19363 14519 19369
rect 14461 19360 14473 19363
rect 14148 19332 14473 19360
rect 14148 19320 14154 19332
rect 14461 19329 14473 19332
rect 14507 19329 14519 19363
rect 14461 19323 14519 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19360 15255 19363
rect 16666 19360 16672 19372
rect 15243 19332 16672 19360
rect 15243 19329 15255 19332
rect 15197 19323 15255 19329
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17218 19320 17224 19372
rect 17276 19320 17282 19372
rect 18892 19369 18920 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 21468 19437 21496 19468
rect 22186 19456 22192 19468
rect 22244 19456 22250 19508
rect 22462 19456 22468 19508
rect 22520 19456 22526 19508
rect 23753 19499 23811 19505
rect 23753 19465 23765 19499
rect 23799 19496 23811 19499
rect 23934 19496 23940 19508
rect 23799 19468 23940 19496
rect 23799 19465 23811 19468
rect 23753 19459 23811 19465
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 25225 19499 25283 19505
rect 25225 19496 25237 19499
rect 24044 19468 25237 19496
rect 21453 19431 21511 19437
rect 21453 19397 21465 19431
rect 21499 19397 21511 19431
rect 21453 19391 21511 19397
rect 21634 19388 21640 19440
rect 21692 19428 21698 19440
rect 24044 19428 24072 19468
rect 25225 19465 25237 19468
rect 25271 19496 25283 19499
rect 25314 19496 25320 19508
rect 25271 19468 25320 19496
rect 25271 19465 25283 19468
rect 25225 19459 25283 19465
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 25774 19456 25780 19508
rect 25832 19456 25838 19508
rect 21692 19400 22140 19428
rect 21692 19388 21698 19400
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19242 19360 19248 19372
rect 19107 19332 19248 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19360 21879 19363
rect 21910 19360 21916 19372
rect 21867 19332 21916 19360
rect 21867 19329 21879 19332
rect 21821 19323 21879 19329
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22112 19369 22140 19400
rect 23584 19400 24072 19428
rect 24112 19431 24170 19437
rect 23584 19369 23612 19400
rect 24112 19397 24124 19431
rect 24158 19428 24170 19431
rect 24394 19428 24400 19440
rect 24158 19400 24400 19428
rect 24158 19397 24170 19400
rect 24112 19391 24170 19397
rect 24394 19388 24400 19400
rect 24452 19388 24458 19440
rect 24854 19388 24860 19440
rect 24912 19428 24918 19440
rect 24912 19400 25636 19428
rect 24912 19388 24918 19400
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19329 23627 19363
rect 23569 19323 23627 19329
rect 5920 19264 6776 19292
rect 8478 19252 8484 19304
rect 8536 19252 8542 19304
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8720 19264 8861 19292
rect 8720 19252 8726 19264
rect 8849 19261 8861 19264
rect 8895 19261 8907 19295
rect 8849 19255 8907 19261
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 7466 19224 7472 19236
rect 5644 19196 7472 19224
rect 4203 19193 4215 19196
rect 4157 19187 4215 19193
rect 7466 19184 7472 19196
rect 7524 19224 7530 19236
rect 7926 19224 7932 19236
rect 7524 19196 7932 19224
rect 7524 19184 7530 19196
rect 7926 19184 7932 19196
rect 7984 19224 7990 19236
rect 8110 19224 8116 19236
rect 7984 19196 8116 19224
rect 7984 19184 7990 19196
rect 8110 19184 8116 19196
rect 8168 19224 8174 19236
rect 10410 19224 10416 19236
rect 8168 19196 10416 19224
rect 8168 19184 8174 19196
rect 10410 19184 10416 19196
rect 10468 19184 10474 19236
rect 2590 19116 2596 19168
rect 2648 19116 2654 19168
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 4798 19156 4804 19168
rect 4755 19128 4804 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 4798 19116 4804 19128
rect 4856 19156 4862 19168
rect 5537 19159 5595 19165
rect 5537 19156 5549 19159
rect 4856 19128 5549 19156
rect 4856 19116 4862 19128
rect 5537 19125 5549 19128
rect 5583 19125 5595 19159
rect 5537 19119 5595 19125
rect 5905 19159 5963 19165
rect 5905 19125 5917 19159
rect 5951 19156 5963 19159
rect 5994 19156 6000 19168
rect 5951 19128 6000 19156
rect 5951 19125 5963 19128
rect 5905 19119 5963 19125
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 7006 19116 7012 19168
rect 7064 19116 7070 19168
rect 8757 19159 8815 19165
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 10318 19156 10324 19168
rect 8803 19128 10324 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10778 19116 10784 19168
rect 10836 19116 10842 19168
rect 10980 19156 11008 19255
rect 13262 19252 13268 19304
rect 13320 19252 13326 19304
rect 13630 19252 13636 19304
rect 13688 19292 13694 19304
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 13688 19264 14565 19292
rect 13688 19252 13694 19264
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14553 19255 14611 19261
rect 15286 19252 15292 19304
rect 15344 19252 15350 19304
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 15654 19252 15660 19304
rect 15712 19292 15718 19304
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 15712 19264 17969 19292
rect 15712 19252 15718 19264
rect 17957 19261 17969 19264
rect 18003 19292 18015 19295
rect 18046 19292 18052 19304
rect 18003 19264 18052 19292
rect 18003 19261 18015 19264
rect 17957 19255 18015 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 22020 19292 22048 19323
rect 22020 19264 22094 19292
rect 22066 19236 22094 19264
rect 13814 19224 13820 19236
rect 12820 19196 13820 19224
rect 12820 19156 12848 19196
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 22066 19196 22100 19236
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 10980 19128 12848 19156
rect 13998 19116 14004 19168
rect 14056 19116 14062 19168
rect 21082 19116 21088 19168
rect 21140 19116 21146 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21269 19159 21327 19165
rect 21269 19156 21281 19159
rect 21232 19128 21281 19156
rect 21232 19116 21238 19128
rect 21269 19125 21281 19128
rect 21315 19125 21327 19159
rect 21269 19119 21327 19125
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 22002 19156 22008 19168
rect 21600 19128 22008 19156
rect 21600 19116 21606 19128
rect 22002 19116 22008 19128
rect 22060 19156 22066 19168
rect 22204 19156 22232 19323
rect 23750 19320 23756 19372
rect 23808 19360 23814 19372
rect 23845 19363 23903 19369
rect 23845 19360 23857 19363
rect 23808 19332 23857 19360
rect 23808 19320 23814 19332
rect 23845 19329 23857 19332
rect 23891 19329 23903 19363
rect 23845 19323 23903 19329
rect 25498 19320 25504 19372
rect 25556 19320 25562 19372
rect 25608 19369 25636 19400
rect 25593 19363 25651 19369
rect 25593 19329 25605 19363
rect 25639 19329 25651 19363
rect 25593 19323 25651 19329
rect 22554 19156 22560 19168
rect 22060 19128 22560 19156
rect 22060 19116 22066 19128
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 25314 19116 25320 19168
rect 25372 19116 25378 19168
rect 1104 19066 26220 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 26220 19066
rect 1104 18992 26220 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 4154 18952 4160 18964
rect 1627 18924 4160 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 5132 18924 5457 18952
rect 5132 18912 5138 18924
rect 5445 18921 5457 18924
rect 5491 18921 5503 18955
rect 10502 18952 10508 18964
rect 5445 18915 5503 18921
rect 5549 18924 10508 18952
rect 2682 18844 2688 18896
rect 2740 18884 2746 18896
rect 5549 18884 5577 18924
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 11701 18955 11759 18961
rect 11701 18921 11713 18955
rect 11747 18952 11759 18955
rect 12253 18955 12311 18961
rect 12253 18952 12265 18955
rect 11747 18924 12265 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 12253 18921 12265 18924
rect 12299 18952 12311 18955
rect 12526 18952 12532 18964
rect 12299 18924 12532 18952
rect 12299 18921 12311 18924
rect 12253 18915 12311 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 13814 18912 13820 18964
rect 13872 18912 13878 18964
rect 16666 18912 16672 18964
rect 16724 18912 16730 18964
rect 21545 18955 21603 18961
rect 21545 18921 21557 18955
rect 21591 18952 21603 18955
rect 22462 18952 22468 18964
rect 21591 18924 22468 18952
rect 21591 18921 21603 18924
rect 21545 18915 21603 18921
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 23661 18955 23719 18961
rect 23661 18921 23673 18955
rect 23707 18952 23719 18955
rect 24486 18952 24492 18964
rect 23707 18924 24492 18952
rect 23707 18921 23719 18924
rect 23661 18915 23719 18921
rect 24486 18912 24492 18924
rect 24544 18912 24550 18964
rect 2740 18856 5577 18884
rect 2740 18844 2746 18856
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 2498 18816 2504 18828
rect 2271 18788 2504 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 2590 18776 2596 18828
rect 2648 18816 2654 18828
rect 3028 18819 3086 18825
rect 3028 18816 3040 18819
rect 2648 18788 3040 18816
rect 2648 18776 2654 18788
rect 3028 18785 3040 18788
rect 3074 18785 3086 18819
rect 3028 18779 3086 18785
rect 3142 18776 3148 18828
rect 3200 18776 3206 18828
rect 3528 18825 3556 18856
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 8478 18884 8484 18896
rect 7892 18856 8484 18884
rect 7892 18844 7898 18856
rect 8478 18844 8484 18856
rect 8536 18884 8542 18896
rect 8536 18856 8616 18884
rect 8536 18844 8542 18856
rect 3513 18819 3571 18825
rect 3513 18785 3525 18819
rect 3559 18785 3571 18819
rect 3513 18779 3571 18785
rect 5626 18776 5632 18828
rect 5684 18776 5690 18828
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 6730 18816 6736 18828
rect 5776 18788 6736 18816
rect 5776 18776 5782 18788
rect 842 18708 848 18760
rect 900 18748 906 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 900 18720 1409 18748
rect 900 18708 906 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2314 18748 2320 18760
rect 2179 18720 2320 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 2516 18748 2544 18776
rect 3237 18751 3295 18757
rect 3237 18748 3249 18751
rect 2516 18720 3249 18748
rect 3237 18717 3249 18720
rect 3283 18717 3295 18751
rect 3237 18711 3295 18717
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 3881 18751 3939 18757
rect 3881 18748 3893 18751
rect 3844 18720 3893 18748
rect 3844 18708 3850 18720
rect 3881 18717 3893 18720
rect 3927 18717 3939 18751
rect 3881 18711 3939 18717
rect 4062 18708 4068 18760
rect 4120 18708 4126 18760
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4798 18708 4804 18760
rect 4856 18708 4862 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18717 5043 18751
rect 4985 18711 5043 18717
rect 2685 18683 2743 18689
rect 2685 18649 2697 18683
rect 2731 18680 2743 18683
rect 2774 18680 2780 18692
rect 2731 18652 2780 18680
rect 2731 18649 2743 18652
rect 2685 18643 2743 18649
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 5000 18680 5028 18711
rect 5074 18708 5080 18760
rect 5132 18708 5138 18760
rect 5350 18757 5356 18760
rect 5341 18751 5356 18757
rect 5341 18717 5353 18751
rect 5341 18711 5356 18717
rect 5350 18708 5356 18711
rect 5408 18708 5414 18760
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6546 18748 6552 18760
rect 5920 18720 6552 18748
rect 5534 18680 5540 18692
rect 5000 18652 5540 18680
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 5920 18680 5948 18720
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 6656 18757 6684 18788
rect 6730 18776 6736 18788
rect 6788 18816 6794 18828
rect 6788 18788 8064 18816
rect 6788 18776 6794 18788
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 8036 18757 8064 18788
rect 8386 18776 8392 18828
rect 8444 18776 8450 18828
rect 8588 18825 8616 18856
rect 10778 18844 10784 18896
rect 10836 18884 10842 18896
rect 12434 18884 12440 18896
rect 10836 18856 12440 18884
rect 10836 18844 10842 18856
rect 12434 18844 12440 18856
rect 12492 18844 12498 18896
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18785 8631 18819
rect 8573 18779 8631 18785
rect 12342 18776 12348 18828
rect 12400 18816 12406 18828
rect 12544 18816 12572 18912
rect 13265 18887 13323 18893
rect 13265 18853 13277 18887
rect 13311 18853 13323 18887
rect 13265 18847 13323 18853
rect 12400 18776 12434 18816
rect 12544 18788 12940 18816
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 7432 18720 7757 18748
rect 7432 18708 7438 18720
rect 7745 18717 7757 18720
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 8021 18751 8079 18757
rect 8021 18717 8033 18751
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 8938 18748 8944 18760
rect 8527 18720 8944 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 5828 18652 5948 18680
rect 1946 18572 1952 18624
rect 2004 18572 2010 18624
rect 2866 18572 2872 18624
rect 2924 18572 2930 18624
rect 3973 18615 4031 18621
rect 3973 18581 3985 18615
rect 4019 18612 4031 18615
rect 4430 18612 4436 18624
rect 4019 18584 4436 18612
rect 4019 18581 4031 18584
rect 3973 18575 4031 18581
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5828 18612 5856 18652
rect 6454 18640 6460 18692
rect 6512 18640 6518 18692
rect 8312 18680 8340 18711
rect 8938 18708 8944 18720
rect 8996 18708 9002 18760
rect 10226 18708 10232 18760
rect 10284 18748 10290 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 10284 18720 10333 18748
rect 10284 18708 10290 18720
rect 10321 18717 10333 18720
rect 10367 18717 10379 18751
rect 12406 18748 12434 18776
rect 12912 18757 12940 18788
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 10321 18711 10379 18717
rect 12084 18720 12817 18748
rect 12084 18692 12112 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 12989 18751 13047 18757
rect 12989 18717 13001 18751
rect 13035 18748 13047 18751
rect 13078 18748 13084 18760
rect 13035 18720 13084 18748
rect 13035 18717 13047 18720
rect 12989 18711 13047 18717
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 13280 18748 13308 18847
rect 22554 18844 22560 18896
rect 22612 18884 22618 18896
rect 22612 18856 22784 18884
rect 22612 18844 22618 18856
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13412 18788 13553 18816
rect 13412 18776 13418 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 15194 18776 15200 18828
rect 15252 18776 15258 18828
rect 17126 18776 17132 18828
rect 17184 18776 17190 18828
rect 17310 18776 17316 18828
rect 17368 18776 17374 18828
rect 22002 18776 22008 18828
rect 22060 18816 22066 18828
rect 22060 18788 22692 18816
rect 22060 18776 22066 18788
rect 13219 18720 13308 18748
rect 13449 18751 13507 18757
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 7484 18652 8984 18680
rect 5307 18584 5856 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 5997 18615 6055 18621
rect 5997 18612 6009 18615
rect 5960 18584 6009 18612
rect 5960 18572 5966 18584
rect 5997 18581 6009 18584
rect 6043 18581 6055 18615
rect 5997 18575 6055 18581
rect 6270 18572 6276 18624
rect 6328 18572 6334 18624
rect 6472 18612 6500 18640
rect 7484 18612 7512 18652
rect 6472 18584 7512 18612
rect 7558 18572 7564 18624
rect 7616 18572 7622 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8386 18612 8392 18624
rect 7975 18584 8392 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 8754 18572 8760 18624
rect 8812 18572 8818 18624
rect 8956 18621 8984 18652
rect 9674 18640 9680 18692
rect 9732 18680 9738 18692
rect 10054 18683 10112 18689
rect 10054 18680 10066 18683
rect 9732 18652 10066 18680
rect 9732 18640 9738 18652
rect 10054 18649 10066 18652
rect 10100 18649 10112 18683
rect 10054 18643 10112 18649
rect 11517 18683 11575 18689
rect 11517 18649 11529 18683
rect 11563 18680 11575 18683
rect 12066 18680 12072 18692
rect 11563 18652 12072 18680
rect 11563 18649 11575 18652
rect 11517 18643 11575 18649
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 12250 18640 12256 18692
rect 12308 18689 12314 18692
rect 12308 18683 12327 18689
rect 12315 18649 12327 18683
rect 13464 18680 13492 18711
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 13909 18751 13967 18757
rect 13909 18748 13921 18751
rect 13688 18720 13921 18748
rect 13688 18708 13694 18720
rect 13909 18717 13921 18720
rect 13955 18717 13967 18751
rect 13909 18711 13967 18717
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14458 18748 14464 18760
rect 14415 18720 14464 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 14608 18720 15853 18748
rect 14608 18708 14614 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 16908 18720 17785 18748
rect 16908 18708 16914 18720
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 20772 18720 21189 18748
rect 20772 18708 20778 18720
rect 21177 18717 21189 18720
rect 21223 18717 21235 18751
rect 21177 18711 21235 18717
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18748 21419 18751
rect 21450 18748 21456 18760
rect 21407 18720 21456 18748
rect 21407 18717 21419 18720
rect 21361 18711 21419 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21542 18708 21548 18760
rect 21600 18748 21606 18760
rect 21821 18751 21879 18757
rect 21600 18747 21772 18748
rect 21821 18747 21833 18751
rect 21600 18720 21833 18747
rect 21600 18708 21606 18720
rect 21744 18719 21833 18720
rect 21821 18717 21833 18719
rect 21867 18717 21879 18751
rect 21821 18711 21879 18717
rect 21913 18729 21971 18735
rect 21913 18695 21925 18729
rect 21959 18695 21971 18729
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 22664 18757 22692 18788
rect 22756 18757 22784 18856
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 24949 18819 25007 18825
rect 24949 18816 24961 18819
rect 23624 18788 24961 18816
rect 23624 18776 23630 18788
rect 24949 18785 24961 18788
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 22557 18751 22615 18757
rect 22557 18748 22569 18751
rect 22480 18720 22569 18748
rect 12308 18643 12327 18649
rect 12452 18652 13492 18680
rect 15381 18683 15439 18689
rect 12308 18640 12314 18643
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 11698 18572 11704 18624
rect 11756 18621 11762 18624
rect 11756 18615 11775 18621
rect 11763 18581 11775 18615
rect 11756 18575 11775 18581
rect 11756 18572 11762 18575
rect 11882 18572 11888 18624
rect 11940 18572 11946 18624
rect 12452 18621 12480 18652
rect 15381 18649 15393 18683
rect 15427 18680 15439 18683
rect 17862 18680 17868 18692
rect 15427 18652 17868 18680
rect 15427 18649 15439 18652
rect 15381 18643 15439 18649
rect 17862 18640 17868 18652
rect 17920 18640 17926 18692
rect 21913 18689 21971 18695
rect 12437 18615 12495 18621
rect 12437 18581 12449 18615
rect 12483 18581 12495 18615
rect 12437 18575 12495 18581
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12986 18612 12992 18624
rect 12575 18584 12992 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 14921 18615 14979 18621
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15289 18615 15347 18621
rect 15289 18612 15301 18615
rect 14967 18584 15301 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15289 18581 15301 18584
rect 15335 18581 15347 18615
rect 15289 18575 15347 18581
rect 15562 18572 15568 18624
rect 15620 18612 15626 18624
rect 15749 18615 15807 18621
rect 15749 18612 15761 18615
rect 15620 18584 15761 18612
rect 15620 18572 15626 18584
rect 15749 18581 15761 18584
rect 15795 18581 15807 18615
rect 15749 18575 15807 18581
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16485 18615 16543 18621
rect 16485 18612 16497 18615
rect 16080 18584 16497 18612
rect 16080 18572 16086 18584
rect 16485 18581 16497 18584
rect 16531 18581 16543 18615
rect 16485 18575 16543 18581
rect 17037 18615 17095 18621
rect 17037 18581 17049 18615
rect 17083 18612 17095 18615
rect 17126 18612 17132 18624
rect 17083 18584 17132 18612
rect 17083 18581 17095 18584
rect 17037 18575 17095 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 18598 18612 18604 18624
rect 18463 18584 18604 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 19610 18572 19616 18624
rect 19668 18612 19674 18624
rect 20254 18612 20260 18624
rect 19668 18584 20260 18612
rect 19668 18572 19674 18584
rect 20254 18572 20260 18584
rect 20312 18612 20318 18624
rect 21358 18612 21364 18624
rect 20312 18584 21364 18612
rect 20312 18572 20318 18584
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 21634 18572 21640 18624
rect 21692 18572 21698 18624
rect 21818 18572 21824 18624
rect 21876 18612 21882 18624
rect 21928 18612 21956 18689
rect 22186 18640 22192 18692
rect 22244 18640 22250 18692
rect 21876 18584 21956 18612
rect 21876 18572 21882 18584
rect 22002 18572 22008 18624
rect 22060 18612 22066 18624
rect 22480 18612 22508 18720
rect 22557 18717 22569 18720
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 22649 18751 22707 18757
rect 22649 18717 22661 18751
rect 22695 18717 22707 18751
rect 22649 18711 22707 18717
rect 22741 18751 22799 18757
rect 22741 18717 22753 18751
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18748 23167 18751
rect 23198 18748 23204 18760
rect 23155 18720 23204 18748
rect 23155 18717 23167 18720
rect 23109 18711 23167 18717
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18748 23535 18751
rect 23658 18748 23664 18760
rect 23523 18720 23664 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 25130 18708 25136 18760
rect 25188 18748 25194 18760
rect 25498 18748 25504 18760
rect 25188 18720 25504 18748
rect 25188 18708 25194 18720
rect 25498 18708 25504 18720
rect 25556 18748 25562 18760
rect 25777 18751 25835 18757
rect 25777 18748 25789 18751
rect 25556 18720 25789 18748
rect 25556 18708 25562 18720
rect 25777 18717 25789 18720
rect 25823 18717 25835 18751
rect 25777 18711 25835 18717
rect 22922 18640 22928 18692
rect 22980 18680 22986 18692
rect 23293 18683 23351 18689
rect 23293 18680 23305 18683
rect 22980 18652 23305 18680
rect 22980 18640 22986 18652
rect 23293 18649 23305 18652
rect 23339 18649 23351 18683
rect 23293 18643 23351 18649
rect 23385 18683 23443 18689
rect 23385 18649 23397 18683
rect 23431 18680 23443 18683
rect 24210 18680 24216 18692
rect 23431 18652 24216 18680
rect 23431 18649 23443 18652
rect 23385 18643 23443 18649
rect 24210 18640 24216 18652
rect 24268 18640 24274 18692
rect 24765 18683 24823 18689
rect 24765 18649 24777 18683
rect 24811 18680 24823 18683
rect 25225 18683 25283 18689
rect 25225 18680 25237 18683
rect 24811 18652 25237 18680
rect 24811 18649 24823 18652
rect 24765 18643 24823 18649
rect 25225 18649 25237 18652
rect 25271 18649 25283 18683
rect 25225 18643 25283 18649
rect 22060 18584 22508 18612
rect 23017 18615 23075 18621
rect 22060 18572 22066 18584
rect 23017 18581 23029 18615
rect 23063 18612 23075 18615
rect 24302 18612 24308 18624
rect 23063 18584 24308 18612
rect 23063 18581 23075 18584
rect 23017 18575 23075 18581
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 24394 18572 24400 18624
rect 24452 18572 24458 18624
rect 24578 18572 24584 18624
rect 24636 18612 24642 18624
rect 24857 18615 24915 18621
rect 24857 18612 24869 18615
rect 24636 18584 24869 18612
rect 24636 18572 24642 18584
rect 24857 18581 24869 18584
rect 24903 18581 24915 18615
rect 24857 18575 24915 18581
rect 1104 18522 26220 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 26220 18522
rect 1104 18448 26220 18470
rect 1857 18411 1915 18417
rect 1857 18377 1869 18411
rect 1903 18408 1915 18411
rect 2222 18408 2228 18420
rect 1903 18380 2228 18408
rect 1903 18377 1915 18380
rect 1857 18371 1915 18377
rect 2222 18368 2228 18380
rect 2280 18408 2286 18420
rect 4062 18408 4068 18420
rect 2280 18380 4068 18408
rect 2280 18368 2286 18380
rect 4062 18368 4068 18380
rect 4120 18408 4126 18420
rect 4985 18411 5043 18417
rect 4120 18380 4752 18408
rect 4120 18368 4126 18380
rect 4724 18349 4752 18380
rect 4985 18377 4997 18411
rect 5031 18408 5043 18411
rect 5258 18408 5264 18420
rect 5031 18380 5264 18408
rect 5031 18377 5043 18380
rect 4985 18371 5043 18377
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5534 18368 5540 18420
rect 5592 18408 5598 18420
rect 7374 18408 7380 18420
rect 5592 18380 7380 18408
rect 5592 18368 5598 18380
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 8168 18380 8309 18408
rect 8168 18368 8174 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 8444 18380 8677 18408
rect 8444 18368 8450 18380
rect 8665 18377 8677 18380
rect 8711 18377 8723 18411
rect 8665 18371 8723 18377
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 8904 18380 10517 18408
rect 8904 18368 8910 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 12250 18368 12256 18420
rect 12308 18408 12314 18420
rect 12345 18411 12403 18417
rect 12345 18408 12357 18411
rect 12308 18380 12357 18408
rect 12308 18368 12314 18380
rect 12345 18377 12357 18380
rect 12391 18377 12403 18411
rect 12345 18371 12403 18377
rect 12434 18368 12440 18420
rect 12492 18368 12498 18420
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 13078 18408 13084 18420
rect 12943 18380 13084 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13538 18368 13544 18420
rect 13596 18368 13602 18420
rect 13814 18368 13820 18420
rect 13872 18368 13878 18420
rect 14001 18411 14059 18417
rect 14001 18377 14013 18411
rect 14047 18408 14059 18411
rect 14458 18408 14464 18420
rect 14047 18380 14464 18408
rect 14047 18377 14059 18380
rect 14001 18371 14059 18377
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19392 18380 19809 18408
rect 19392 18368 19398 18380
rect 19797 18377 19809 18380
rect 19843 18408 19855 18411
rect 20622 18408 20628 18420
rect 19843 18380 20628 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 20622 18368 20628 18380
rect 20680 18408 20686 18420
rect 21818 18408 21824 18420
rect 20680 18380 21824 18408
rect 20680 18368 20686 18380
rect 21818 18368 21824 18380
rect 21876 18368 21882 18420
rect 23198 18368 23204 18420
rect 23256 18408 23262 18420
rect 23293 18411 23351 18417
rect 23293 18408 23305 18411
rect 23256 18380 23305 18408
rect 23256 18368 23262 18380
rect 23293 18377 23305 18380
rect 23339 18377 23351 18411
rect 23293 18371 23351 18377
rect 25130 18368 25136 18420
rect 25188 18368 25194 18420
rect 25406 18368 25412 18420
rect 25464 18368 25470 18420
rect 4341 18343 4399 18349
rect 2746 18312 3280 18340
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 2746 18272 2774 18312
rect 2464 18244 2774 18272
rect 2464 18232 2470 18244
rect 2958 18232 2964 18284
rect 3016 18281 3022 18284
rect 3252 18281 3280 18312
rect 4341 18309 4353 18343
rect 4387 18340 4399 18343
rect 4617 18343 4675 18349
rect 4617 18340 4629 18343
rect 4387 18312 4629 18340
rect 4387 18309 4399 18312
rect 4341 18303 4399 18309
rect 4617 18309 4629 18312
rect 4663 18309 4675 18343
rect 4617 18303 4675 18309
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18309 4767 18343
rect 5718 18340 5724 18352
rect 4709 18303 4767 18309
rect 4816 18312 5724 18340
rect 3016 18272 3028 18281
rect 3237 18275 3295 18281
rect 3016 18244 3061 18272
rect 3016 18235 3028 18244
rect 3237 18241 3249 18275
rect 3283 18241 3295 18275
rect 3237 18235 3295 18241
rect 3016 18232 3022 18235
rect 3970 18232 3976 18284
rect 4028 18232 4034 18284
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4120 18244 4165 18272
rect 4120 18232 4126 18244
rect 4430 18232 4436 18284
rect 4488 18232 4494 18284
rect 4816 18281 4844 18312
rect 5718 18300 5724 18312
rect 5776 18300 5782 18352
rect 6454 18340 6460 18352
rect 5828 18312 6460 18340
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18241 4859 18275
rect 4801 18235 4859 18241
rect 5534 18275 5592 18281
rect 5534 18241 5546 18275
rect 5580 18272 5592 18275
rect 5828 18272 5856 18312
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 7926 18340 7932 18352
rect 7340 18312 7932 18340
rect 7340 18300 7346 18312
rect 5580 18244 5856 18272
rect 5580 18241 5592 18244
rect 5534 18235 5592 18241
rect 5902 18232 5908 18284
rect 5960 18232 5966 18284
rect 5994 18232 6000 18284
rect 6052 18232 6058 18284
rect 6914 18232 6920 18284
rect 6972 18232 6978 18284
rect 7190 18232 7196 18284
rect 7248 18232 7254 18284
rect 7668 18281 7696 18312
rect 7926 18300 7932 18312
rect 7984 18340 7990 18352
rect 8404 18340 8432 18368
rect 10318 18349 10324 18352
rect 7984 18312 8432 18340
rect 10296 18343 10324 18349
rect 7984 18300 7990 18312
rect 10296 18309 10308 18343
rect 10296 18303 10324 18309
rect 10318 18300 10324 18303
rect 10376 18300 10382 18352
rect 10410 18300 10416 18352
rect 10468 18300 10474 18352
rect 12452 18340 12480 18368
rect 13446 18340 13452 18352
rect 12452 18312 13452 18340
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18204 6791 18207
rect 7006 18204 7012 18216
rect 6779 18176 7012 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7484 18204 7512 18235
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 8414 18275 8472 18281
rect 8414 18241 8426 18275
rect 8460 18272 8472 18275
rect 8570 18272 8576 18284
rect 8460 18244 8576 18272
rect 8460 18241 8472 18244
rect 8414 18235 8472 18241
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 9789 18275 9847 18281
rect 9789 18241 9801 18275
rect 9835 18272 9847 18275
rect 9835 18244 10272 18272
rect 9835 18241 9847 18244
rect 9789 18235 9847 18241
rect 7156 18176 7512 18204
rect 7156 18164 7162 18176
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 7929 18207 7987 18213
rect 7929 18204 7941 18207
rect 7800 18176 7941 18204
rect 7800 18164 7806 18176
rect 7929 18173 7941 18176
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 8202 18164 8208 18216
rect 8260 18164 8266 18216
rect 10045 18207 10103 18213
rect 10045 18173 10057 18207
rect 10091 18204 10103 18207
rect 10134 18204 10140 18216
rect 10091 18176 10140 18204
rect 10091 18173 10103 18176
rect 10045 18167 10103 18173
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 7285 18139 7343 18145
rect 7285 18105 7297 18139
rect 7331 18136 7343 18139
rect 8220 18136 8248 18164
rect 7331 18108 8248 18136
rect 8573 18139 8631 18145
rect 7331 18105 7343 18108
rect 7285 18099 7343 18105
rect 8573 18105 8585 18139
rect 8619 18136 8631 18139
rect 10244 18136 10272 18244
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12308 18244 12449 18272
rect 12308 18232 12314 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10560 18176 10793 18204
rect 10560 18164 10566 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12342 18204 12348 18216
rect 11931 18176 12348 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12342 18164 12348 18176
rect 12400 18164 12406 18216
rect 12618 18164 12624 18216
rect 12676 18164 12682 18216
rect 12728 18204 12756 18235
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 13096 18281 13124 18312
rect 13446 18300 13452 18312
rect 13504 18300 13510 18352
rect 15562 18300 15568 18352
rect 15620 18349 15626 18352
rect 15620 18340 15632 18349
rect 17988 18343 18046 18349
rect 15620 18312 15665 18340
rect 15620 18303 15632 18312
rect 17988 18309 18000 18343
rect 18034 18340 18046 18343
rect 18325 18343 18383 18349
rect 18325 18340 18337 18343
rect 18034 18312 18337 18340
rect 18034 18309 18046 18312
rect 17988 18303 18046 18309
rect 18325 18309 18337 18312
rect 18371 18309 18383 18343
rect 20257 18343 20315 18349
rect 20257 18340 20269 18343
rect 18325 18303 18383 18309
rect 18800 18312 20269 18340
rect 15620 18300 15626 18303
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 13170 18232 13176 18284
rect 13228 18272 13234 18284
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 13228 18244 13277 18272
rect 13228 18232 13234 18244
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 13998 18272 14004 18284
rect 13403 18244 14004 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14366 18232 14372 18284
rect 14424 18232 14430 18284
rect 15746 18232 15752 18284
rect 15804 18272 15810 18284
rect 15841 18275 15899 18281
rect 15841 18272 15853 18275
rect 15804 18244 15853 18272
rect 15804 18232 15810 18244
rect 15841 18241 15853 18244
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18196 18244 18245 18272
rect 18196 18232 18202 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 13630 18204 13636 18216
rect 12728 18176 13636 18204
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 18524 18204 18552 18235
rect 18598 18232 18604 18284
rect 18656 18232 18662 18284
rect 18800 18213 18828 18312
rect 20257 18309 20269 18312
rect 20303 18340 20315 18343
rect 23109 18343 23167 18349
rect 20303 18312 22048 18340
rect 20303 18309 20315 18312
rect 20257 18303 20315 18309
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18272 18935 18275
rect 19058 18272 19064 18284
rect 18923 18244 19064 18272
rect 18923 18241 18935 18244
rect 18877 18235 18935 18241
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 19610 18232 19616 18284
rect 19668 18232 19674 18284
rect 19886 18232 19892 18284
rect 19944 18272 19950 18284
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 19944 18244 20085 18272
rect 19944 18232 19950 18244
rect 20073 18241 20085 18244
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 20162 18232 20168 18284
rect 20220 18232 20226 18284
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 18785 18207 18843 18213
rect 18524 18176 18644 18204
rect 8619 18108 9168 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 5353 18071 5411 18077
rect 5353 18037 5365 18071
rect 5399 18068 5411 18071
rect 7466 18068 7472 18080
rect 5399 18040 7472 18068
rect 5399 18037 5411 18040
rect 5353 18031 5411 18037
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18068 7803 18071
rect 8478 18068 8484 18080
rect 7791 18040 8484 18068
rect 7791 18037 7803 18040
rect 7745 18031 7803 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 9140 18068 9168 18108
rect 10152 18108 10272 18136
rect 12253 18139 12311 18145
rect 10042 18068 10048 18080
rect 9140 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10152 18077 10180 18108
rect 12253 18105 12265 18139
rect 12299 18136 12311 18139
rect 12894 18136 12900 18148
rect 12299 18108 12900 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 12894 18096 12900 18108
rect 12952 18096 12958 18148
rect 10137 18071 10195 18077
rect 10137 18037 10149 18071
rect 10183 18037 10195 18071
rect 10137 18031 10195 18037
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 11940 18040 12449 18068
rect 11940 18028 11946 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12437 18031 12495 18037
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 14001 18071 14059 18077
rect 14001 18068 14013 18071
rect 12584 18040 14013 18068
rect 12584 18028 12590 18040
rect 14001 18037 14013 18040
rect 14047 18037 14059 18071
rect 14001 18031 14059 18037
rect 16850 18028 16856 18080
rect 16908 18028 16914 18080
rect 18616 18068 18644 18176
rect 18785 18173 18797 18207
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 19484 18176 19993 18204
rect 19484 18164 19490 18176
rect 19981 18173 19993 18176
rect 20027 18204 20039 18207
rect 20180 18204 20208 18232
rect 20027 18176 20208 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20364 18204 20392 18235
rect 20312 18176 20392 18204
rect 20456 18204 20484 18235
rect 20530 18232 20536 18284
rect 20588 18232 20594 18284
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20640 18204 20668 18235
rect 20714 18232 20720 18284
rect 20772 18232 20778 18284
rect 20898 18232 20904 18284
rect 20956 18232 20962 18284
rect 21450 18272 21456 18284
rect 21100 18244 21456 18272
rect 20809 18207 20867 18213
rect 20809 18204 20821 18207
rect 20456 18176 20576 18204
rect 20640 18176 20821 18204
rect 20312 18164 20318 18176
rect 20070 18096 20076 18148
rect 20128 18136 20134 18148
rect 20548 18136 20576 18176
rect 20809 18173 20821 18176
rect 20855 18204 20867 18207
rect 21100 18204 21128 18244
rect 21450 18232 21456 18244
rect 21508 18272 21514 18284
rect 21545 18275 21603 18281
rect 21545 18272 21557 18275
rect 21508 18244 21557 18272
rect 21508 18232 21514 18244
rect 21545 18241 21557 18244
rect 21591 18241 21603 18275
rect 21545 18235 21603 18241
rect 21634 18232 21640 18284
rect 21692 18232 21698 18284
rect 21818 18232 21824 18284
rect 21876 18232 21882 18284
rect 21913 18275 21971 18281
rect 21913 18241 21925 18275
rect 21959 18241 21971 18275
rect 21913 18235 21971 18241
rect 20855 18176 21128 18204
rect 20855 18173 20867 18176
rect 20809 18167 20867 18173
rect 21174 18164 21180 18216
rect 21232 18164 21238 18216
rect 21928 18204 21956 18235
rect 21836 18176 21956 18204
rect 22020 18204 22048 18312
rect 23109 18309 23121 18343
rect 23155 18340 23167 18343
rect 24020 18343 24078 18349
rect 23155 18312 23796 18340
rect 23155 18309 23167 18312
rect 23109 18303 23167 18309
rect 23768 18284 23796 18312
rect 24020 18309 24032 18343
rect 24066 18340 24078 18343
rect 24394 18340 24400 18352
rect 24066 18312 24400 18340
rect 24066 18309 24078 18312
rect 24020 18303 24078 18309
rect 24394 18300 24400 18312
rect 24452 18300 24458 18352
rect 22278 18232 22284 18284
rect 22336 18232 22342 18284
rect 22738 18232 22744 18284
rect 22796 18272 22802 18284
rect 23293 18275 23351 18281
rect 23293 18272 23305 18275
rect 22796 18244 23305 18272
rect 22796 18232 22802 18244
rect 23293 18241 23305 18244
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18241 23535 18275
rect 23477 18235 23535 18241
rect 23492 18204 23520 18235
rect 23750 18232 23756 18284
rect 23808 18232 23814 18284
rect 25225 18275 25283 18281
rect 25225 18241 25237 18275
rect 25271 18272 25283 18275
rect 25314 18272 25320 18284
rect 25271 18244 25320 18272
rect 25271 18241 25283 18244
rect 25225 18235 25283 18241
rect 25314 18232 25320 18244
rect 25372 18232 25378 18284
rect 25590 18232 25596 18284
rect 25648 18232 25654 18284
rect 22020 18176 23520 18204
rect 20128 18108 21312 18136
rect 20128 18096 20134 18108
rect 21284 18080 21312 18108
rect 21358 18096 21364 18148
rect 21416 18096 21422 18148
rect 21836 18136 21864 18176
rect 21910 18136 21916 18148
rect 21836 18108 21916 18136
rect 21910 18096 21916 18108
rect 21968 18136 21974 18148
rect 22738 18136 22744 18148
rect 21968 18108 22744 18136
rect 21968 18096 21974 18108
rect 22738 18096 22744 18108
rect 22796 18096 22802 18148
rect 20438 18068 20444 18080
rect 18616 18040 20444 18068
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 21266 18028 21272 18080
rect 21324 18068 21330 18080
rect 21634 18068 21640 18080
rect 21324 18040 21640 18068
rect 21324 18028 21330 18040
rect 21634 18028 21640 18040
rect 21692 18068 21698 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21692 18040 21833 18068
rect 21692 18028 21698 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22189 18071 22247 18077
rect 22189 18068 22201 18071
rect 22152 18040 22201 18068
rect 22152 18028 22158 18040
rect 22189 18037 22201 18040
rect 22235 18037 22247 18071
rect 22189 18031 22247 18037
rect 25774 18028 25780 18080
rect 25832 18028 25838 18080
rect 1104 17978 26220 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 26220 17978
rect 1104 17904 26220 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2832 17836 2973 17864
rect 2832 17824 2838 17836
rect 2961 17833 2973 17836
rect 3007 17864 3019 17867
rect 3970 17864 3976 17876
rect 3007 17836 3976 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 5350 17824 5356 17876
rect 5408 17864 5414 17876
rect 5445 17867 5503 17873
rect 5445 17864 5457 17867
rect 5408 17836 5457 17864
rect 5408 17824 5414 17836
rect 5445 17833 5457 17836
rect 5491 17833 5503 17867
rect 6822 17864 6828 17876
rect 5445 17827 5503 17833
rect 5549 17836 6828 17864
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 5549 17796 5577 17836
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 6972 17836 7481 17864
rect 6972 17824 6978 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 8665 17867 8723 17873
rect 8665 17833 8677 17867
rect 8711 17864 8723 17867
rect 9674 17864 9680 17876
rect 8711 17836 9680 17864
rect 8711 17833 8723 17836
rect 8665 17827 8723 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 12526 17864 12532 17876
rect 12483 17836 12532 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12618 17824 12624 17876
rect 12676 17824 12682 17876
rect 13173 17867 13231 17873
rect 13173 17833 13185 17867
rect 13219 17864 13231 17867
rect 13354 17864 13360 17876
rect 13219 17836 13360 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 14090 17824 14096 17876
rect 14148 17824 14154 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15252 17836 16068 17864
rect 15252 17824 15258 17836
rect 4212 17768 5577 17796
rect 6365 17799 6423 17805
rect 4212 17756 4218 17768
rect 6365 17765 6377 17799
rect 6411 17796 6423 17799
rect 7190 17796 7196 17808
rect 6411 17768 7196 17796
rect 6411 17765 6423 17768
rect 6365 17759 6423 17765
rect 7190 17756 7196 17768
rect 7248 17756 7254 17808
rect 7742 17756 7748 17808
rect 7800 17796 7806 17808
rect 7800 17768 8064 17796
rect 7800 17756 7806 17768
rect 6270 17728 6276 17740
rect 5644 17700 6276 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 2314 17660 2320 17672
rect 1627 17632 2320 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 2314 17620 2320 17632
rect 2372 17620 2378 17672
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 5644 17669 5672 17700
rect 6270 17688 6276 17700
rect 6328 17728 6334 17740
rect 7101 17731 7159 17737
rect 6328 17700 6868 17728
rect 6328 17688 6334 17700
rect 5629 17663 5687 17669
rect 4028 17632 4292 17660
rect 4028 17620 4034 17632
rect 1848 17595 1906 17601
rect 1848 17561 1860 17595
rect 1894 17592 1906 17595
rect 1946 17592 1952 17604
rect 1894 17564 1952 17592
rect 1894 17561 1906 17564
rect 1848 17555 1906 17561
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 4154 17552 4160 17604
rect 4212 17552 4218 17604
rect 4264 17592 4292 17632
rect 5629 17629 5641 17663
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 5905 17663 5963 17669
rect 5905 17629 5917 17663
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 5920 17592 5948 17623
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 6840 17660 6868 17700
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7374 17728 7380 17740
rect 7147 17700 7380 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7374 17688 7380 17700
rect 7432 17728 7438 17740
rect 8036 17737 8064 17768
rect 8938 17756 8944 17808
rect 8996 17756 9002 17808
rect 12066 17756 12072 17808
rect 12124 17756 12130 17808
rect 8021 17731 8079 17737
rect 7432 17700 7671 17728
rect 7432 17688 7438 17700
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 6687 17632 6776 17660
rect 6840 17632 7021 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 4264 17564 5948 17592
rect 4065 17527 4123 17533
rect 4065 17493 4077 17527
rect 4111 17524 4123 17527
rect 4430 17524 4436 17536
rect 4111 17496 4436 17524
rect 4111 17493 4123 17496
rect 4065 17487 4123 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 6748 17524 6776 17632
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7009 17623 7067 17629
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7282 17620 7288 17672
rect 7340 17620 7346 17672
rect 7643 17669 7671 17700
rect 8021 17697 8033 17731
rect 8067 17697 8079 17731
rect 8021 17691 8079 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8352 17700 8401 17728
rect 8352 17688 8358 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 8506 17731 8564 17737
rect 8506 17697 8518 17731
rect 8552 17728 8564 17731
rect 8754 17728 8760 17740
rect 8552 17700 8760 17728
rect 8552 17697 8564 17700
rect 8506 17691 8564 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 12544 17728 12572 17824
rect 13081 17799 13139 17805
rect 13081 17765 13093 17799
rect 13127 17765 13139 17799
rect 13081 17759 13139 17765
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 12544 17700 12725 17728
rect 12713 17697 12725 17700
rect 12759 17697 12771 17731
rect 12713 17691 12771 17697
rect 7585 17663 7671 17669
rect 7585 17629 7597 17663
rect 7631 17632 7671 17663
rect 7745 17663 7803 17669
rect 7631 17629 7643 17632
rect 7585 17623 7643 17629
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 7926 17660 7932 17672
rect 7791 17632 7932 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 10042 17620 10048 17672
rect 10100 17669 10106 17672
rect 10100 17660 10112 17669
rect 10100 17632 10145 17660
rect 10100 17623 10112 17632
rect 10100 17620 10106 17623
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 10284 17632 10333 17660
rect 10284 17620 10290 17632
rect 10321 17629 10333 17632
rect 10367 17629 10379 17663
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10321 17623 10379 17629
rect 10980 17632 11805 17660
rect 6825 17595 6883 17601
rect 6825 17561 6837 17595
rect 6871 17592 6883 17595
rect 8297 17595 8355 17601
rect 6871 17564 7604 17592
rect 6871 17561 6883 17564
rect 6825 17555 6883 17561
rect 7576 17536 7604 17564
rect 8297 17561 8309 17595
rect 8343 17592 8355 17595
rect 8662 17592 8668 17604
rect 8343 17564 8668 17592
rect 8343 17561 8355 17564
rect 8297 17555 8355 17561
rect 8662 17552 8668 17564
rect 8720 17552 8726 17604
rect 10336 17592 10364 17623
rect 10980 17604 11008 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 10597 17595 10655 17601
rect 10597 17592 10609 17595
rect 10336 17564 10609 17592
rect 10597 17561 10609 17564
rect 10643 17592 10655 17595
rect 10962 17592 10968 17604
rect 10643 17564 10968 17592
rect 10643 17561 10655 17564
rect 10597 17555 10655 17561
rect 10962 17552 10968 17564
rect 11020 17552 11026 17604
rect 11054 17552 11060 17604
rect 11112 17552 11118 17604
rect 13096 17592 13124 17759
rect 13357 17731 13415 17737
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 14108 17728 14136 17824
rect 16040 17796 16068 17836
rect 17862 17824 17868 17876
rect 17920 17824 17926 17876
rect 19334 17824 19340 17876
rect 19392 17824 19398 17876
rect 19794 17824 19800 17876
rect 19852 17864 19858 17876
rect 20530 17864 20536 17876
rect 19852 17836 20536 17864
rect 19852 17824 19858 17836
rect 20530 17824 20536 17836
rect 20588 17824 20594 17876
rect 20990 17824 20996 17876
rect 21048 17864 21054 17876
rect 21266 17864 21272 17876
rect 21048 17836 21272 17864
rect 21048 17824 21054 17836
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 21545 17867 21603 17873
rect 21545 17833 21557 17867
rect 21591 17864 21603 17867
rect 23566 17864 23572 17876
rect 21591 17836 23572 17864
rect 21591 17833 21603 17836
rect 21545 17827 21603 17833
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 17218 17796 17224 17808
rect 16040 17768 16160 17796
rect 16132 17740 16160 17768
rect 16960 17768 17224 17796
rect 16025 17731 16083 17737
rect 16025 17728 16037 17731
rect 13403 17700 14136 17728
rect 15396 17700 16037 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17660 13967 17663
rect 15396 17660 15424 17700
rect 16025 17697 16037 17700
rect 16071 17697 16083 17731
rect 16025 17691 16083 17697
rect 16114 17688 16120 17740
rect 16172 17688 16178 17740
rect 13955 17632 15424 17660
rect 13955 17629 13967 17632
rect 13909 17623 13967 17629
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16632 17632 16865 17660
rect 16632 17620 16638 17632
rect 16853 17629 16865 17632
rect 16899 17660 16911 17663
rect 16960 17660 16988 17768
rect 17218 17756 17224 17768
rect 17276 17796 17282 17808
rect 22278 17796 22284 17808
rect 17276 17768 22284 17796
rect 17276 17756 17282 17768
rect 22278 17756 22284 17768
rect 22336 17756 22342 17808
rect 18322 17688 18328 17740
rect 18380 17688 18386 17740
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17697 18475 17731
rect 18417 17691 18475 17697
rect 16899 17632 16988 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17862 17660 17868 17672
rect 17368 17632 17868 17660
rect 17368 17620 17374 17632
rect 17862 17620 17868 17632
rect 17920 17660 17926 17672
rect 18432 17660 18460 17691
rect 19518 17688 19524 17740
rect 19576 17688 19582 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20956 17700 21189 17728
rect 20956 17688 20962 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 21634 17728 21640 17740
rect 21177 17691 21235 17697
rect 21284 17700 21640 17728
rect 17920 17632 18460 17660
rect 17920 17620 17926 17632
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19300 17632 19717 17660
rect 19300 17620 19306 17632
rect 19705 17629 19717 17632
rect 19751 17660 19763 17663
rect 20809 17663 20867 17669
rect 19751 17632 20760 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 14550 17592 14556 17604
rect 13096 17564 14556 17592
rect 14550 17552 14556 17564
rect 14608 17552 14614 17604
rect 15228 17595 15286 17601
rect 15228 17561 15240 17595
rect 15274 17592 15286 17595
rect 15274 17564 15608 17592
rect 15274 17561 15286 17564
rect 15228 17555 15286 17561
rect 7190 17524 7196 17536
rect 6748 17496 7196 17524
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7558 17484 7564 17536
rect 7616 17484 7622 17536
rect 7650 17484 7656 17536
rect 7708 17484 7714 17536
rect 12434 17484 12440 17536
rect 12492 17484 12498 17536
rect 15580 17533 15608 17564
rect 17586 17552 17592 17604
rect 17644 17552 17650 17604
rect 15565 17527 15623 17533
rect 15565 17493 15577 17527
rect 15611 17493 15623 17527
rect 15565 17487 15623 17493
rect 15930 17484 15936 17536
rect 15988 17484 15994 17536
rect 18230 17484 18236 17536
rect 18288 17484 18294 17536
rect 19521 17527 19579 17533
rect 19521 17493 19533 17527
rect 19567 17524 19579 17527
rect 19702 17524 19708 17536
rect 19567 17496 19708 17524
rect 19567 17493 19579 17496
rect 19521 17487 19579 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 20732 17524 20760 17632
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 20824 17592 20852 17623
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17662 21143 17663
rect 21284 17662 21312 17700
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 24302 17688 24308 17740
rect 24360 17728 24366 17740
rect 24949 17731 25007 17737
rect 24949 17728 24961 17731
rect 24360 17700 24961 17728
rect 24360 17688 24366 17700
rect 24949 17697 24961 17700
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 21131 17634 21312 17662
rect 21361 17663 21419 17669
rect 21131 17629 21143 17634
rect 21085 17623 21143 17629
rect 21361 17629 21373 17663
rect 21407 17660 21419 17663
rect 21542 17660 21548 17672
rect 21407 17632 21548 17660
rect 21407 17629 21419 17632
rect 21361 17623 21419 17629
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 21726 17620 21732 17672
rect 21784 17660 21790 17672
rect 21821 17663 21879 17669
rect 21821 17660 21833 17663
rect 21784 17632 21833 17660
rect 21784 17620 21790 17632
rect 21821 17629 21833 17632
rect 21867 17629 21879 17663
rect 21821 17623 21879 17629
rect 21910 17620 21916 17672
rect 21968 17620 21974 17672
rect 22281 17663 22339 17669
rect 22281 17629 22293 17663
rect 22327 17660 22339 17663
rect 23750 17660 23756 17672
rect 22327 17632 23756 17660
rect 22327 17629 22339 17632
rect 22281 17623 22339 17629
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 25130 17620 25136 17672
rect 25188 17660 25194 17672
rect 25777 17663 25835 17669
rect 25777 17660 25789 17663
rect 25188 17632 25789 17660
rect 25188 17620 25194 17632
rect 25777 17629 25789 17632
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 21174 17592 21180 17604
rect 20824 17564 21180 17592
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 21266 17552 21272 17604
rect 21324 17592 21330 17604
rect 21637 17595 21695 17601
rect 21637 17592 21649 17595
rect 21324 17564 21649 17592
rect 21324 17552 21330 17564
rect 21637 17561 21649 17564
rect 21683 17561 21695 17595
rect 21928 17592 21956 17620
rect 21637 17555 21695 17561
rect 21744 17564 21956 17592
rect 24765 17595 24823 17601
rect 21744 17524 21772 17564
rect 24765 17561 24777 17595
rect 24811 17592 24823 17595
rect 25225 17595 25283 17601
rect 25225 17592 25237 17595
rect 24811 17564 25237 17592
rect 24811 17561 24823 17564
rect 24765 17555 24823 17561
rect 25225 17561 25237 17564
rect 25271 17561 25283 17595
rect 25225 17555 25283 17561
rect 20732 17496 21772 17524
rect 21910 17484 21916 17536
rect 21968 17484 21974 17536
rect 24026 17484 24032 17536
rect 24084 17524 24090 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 24084 17496 24409 17524
rect 24084 17484 24090 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 24397 17487 24455 17493
rect 24486 17484 24492 17536
rect 24544 17524 24550 17536
rect 24857 17527 24915 17533
rect 24857 17524 24869 17527
rect 24544 17496 24869 17524
rect 24544 17484 24550 17496
rect 24857 17493 24869 17496
rect 24903 17493 24915 17527
rect 24857 17487 24915 17493
rect 1104 17434 26220 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 26220 17434
rect 1104 17360 26220 17382
rect 3786 17320 3792 17332
rect 3160 17292 3792 17320
rect 3160 17193 3188 17292
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 4614 17280 4620 17332
rect 4672 17280 4678 17332
rect 7285 17323 7343 17329
rect 7285 17289 7297 17323
rect 7331 17289 7343 17323
rect 7285 17283 7343 17289
rect 8297 17323 8355 17329
rect 8297 17289 8309 17323
rect 8343 17320 8355 17323
rect 8570 17320 8576 17332
rect 8343 17292 8576 17320
rect 8343 17289 8355 17292
rect 8297 17283 8355 17289
rect 7300 17252 7328 17283
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 14734 17320 14740 17332
rect 11112 17292 14740 17320
rect 11112 17280 11118 17292
rect 14734 17280 14740 17292
rect 14792 17320 14798 17332
rect 16574 17320 16580 17332
rect 14792 17292 16580 17320
rect 14792 17280 14798 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 21082 17320 21088 17332
rect 19628 17292 21088 17320
rect 7377 17255 7435 17261
rect 7377 17252 7389 17255
rect 3252 17224 4446 17252
rect 7300 17224 7389 17252
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 3252 17125 3280 17224
rect 4418 17196 4446 17224
rect 7377 17221 7389 17224
rect 7423 17221 7435 17255
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 7377 17215 7435 17221
rect 7484 17224 7696 17252
rect 3786 17144 3792 17196
rect 3844 17184 3850 17196
rect 4418 17193 4436 17196
rect 4249 17187 4307 17193
rect 4249 17184 4261 17187
rect 3844 17156 4261 17184
rect 3844 17144 3850 17156
rect 4249 17153 4261 17156
rect 4295 17153 4307 17187
rect 4249 17147 4307 17153
rect 4403 17187 4436 17193
rect 4403 17153 4415 17187
rect 4488 17184 4494 17196
rect 6270 17184 6276 17196
rect 4488 17156 6276 17184
rect 4403 17147 4436 17153
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 3513 17119 3571 17125
rect 3513 17085 3525 17119
rect 3559 17116 3571 17119
rect 3878 17116 3884 17128
rect 3559 17088 3884 17116
rect 3559 17085 3571 17088
rect 3513 17079 3571 17085
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4264 17116 4292 17147
rect 4430 17144 4436 17147
rect 4488 17144 4494 17156
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7098 17184 7104 17196
rect 6963 17156 7104 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7098 17144 7104 17156
rect 7156 17144 7162 17196
rect 7190 17144 7196 17196
rect 7248 17184 7254 17196
rect 7484 17184 7512 17224
rect 7248 17156 7512 17184
rect 7248 17144 7254 17156
rect 7558 17144 7564 17196
rect 7616 17144 7622 17196
rect 7668 17193 7696 17224
rect 15856 17224 16865 17252
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 7699 17156 8677 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 8665 17153 8677 17156
rect 8711 17184 8723 17187
rect 8938 17184 8944 17196
rect 8711 17156 8944 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 11790 17193 11796 17196
rect 11784 17147 11796 17193
rect 11790 17144 11796 17147
rect 11848 17144 11854 17196
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 12952 17156 13553 17184
rect 12952 17144 12958 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 15217 17187 15275 17193
rect 15217 17153 15229 17187
rect 15263 17184 15275 17187
rect 15263 17156 15424 17184
rect 15263 17153 15275 17156
rect 15217 17147 15275 17153
rect 6178 17116 6184 17128
rect 4264 17088 6184 17116
rect 6178 17076 6184 17088
rect 6236 17116 6242 17128
rect 6380 17116 6408 17144
rect 6236 17088 6408 17116
rect 7009 17119 7067 17125
rect 6236 17076 6242 17088
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7926 17116 7932 17128
rect 7055 17088 7932 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7926 17076 7932 17088
rect 7984 17076 7990 17128
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8573 17119 8631 17125
rect 8573 17116 8585 17119
rect 8536 17088 8585 17116
rect 8536 17076 8542 17088
rect 8573 17085 8585 17088
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11020 17088 11529 17116
rect 11020 17076 11026 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 15396 17116 15424 17156
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15856 17184 15884 17224
rect 16853 17221 16865 17224
rect 16899 17252 16911 17255
rect 16942 17252 16948 17264
rect 16899 17224 16948 17252
rect 16899 17221 16911 17224
rect 16853 17215 16911 17221
rect 16942 17212 16948 17224
rect 17000 17252 17006 17264
rect 17586 17252 17592 17264
rect 17000 17224 17592 17252
rect 17000 17212 17006 17224
rect 17586 17212 17592 17224
rect 17644 17212 17650 17264
rect 18233 17255 18291 17261
rect 18233 17221 18245 17255
rect 18279 17252 18291 17255
rect 18414 17252 18420 17264
rect 18279 17224 18420 17252
rect 18279 17221 18291 17224
rect 18233 17215 18291 17221
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 19153 17255 19211 17261
rect 19153 17221 19165 17255
rect 19199 17252 19211 17255
rect 19426 17252 19432 17264
rect 19199 17224 19432 17252
rect 19199 17221 19211 17224
rect 19153 17215 19211 17221
rect 19426 17212 19432 17224
rect 19484 17212 19490 17264
rect 15528 17156 15884 17184
rect 15933 17187 15991 17193
rect 15528 17144 15534 17156
rect 15933 17153 15945 17187
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 15396 17088 15608 17116
rect 11517 17079 11575 17085
rect 5902 17008 5908 17060
rect 5960 17048 5966 17060
rect 15580 17057 15608 17088
rect 7837 17051 7895 17057
rect 7837 17048 7849 17051
rect 5960 17020 7849 17048
rect 5960 17008 5966 17020
rect 7837 17017 7849 17020
rect 7883 17017 7895 17051
rect 12989 17051 13047 17057
rect 12989 17048 13001 17051
rect 7837 17011 7895 17017
rect 12728 17020 13001 17048
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16980 6515 16983
rect 6546 16980 6552 16992
rect 6503 16952 6552 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 6546 16940 6552 16952
rect 6604 16980 6610 16992
rect 6822 16980 6828 16992
rect 6604 16952 6828 16980
rect 6604 16940 6610 16952
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7650 16940 7656 16992
rect 7708 16940 7714 16992
rect 12250 16940 12256 16992
rect 12308 16980 12314 16992
rect 12728 16980 12756 17020
rect 12989 17017 13001 17020
rect 13035 17017 13047 17051
rect 12989 17011 13047 17017
rect 15565 17051 15623 17057
rect 15565 17017 15577 17051
rect 15611 17017 15623 17051
rect 15948 17048 15976 17147
rect 16022 17144 16028 17196
rect 16080 17144 16086 17196
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 19061 17187 19119 17193
rect 17920 17156 18460 17184
rect 17920 17144 17926 17156
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 18322 17076 18328 17128
rect 18380 17076 18386 17128
rect 18432 17125 18460 17156
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 19107 17156 19533 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19521 17153 19533 17156
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17116 19303 17119
rect 19628 17116 19656 17292
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 22094 17320 22100 17332
rect 21416 17292 22100 17320
rect 21416 17280 21422 17292
rect 22094 17280 22100 17292
rect 22152 17280 22158 17332
rect 22189 17323 22247 17329
rect 22189 17289 22201 17323
rect 22235 17320 22247 17323
rect 22370 17320 22376 17332
rect 22235 17292 22376 17320
rect 22235 17289 22247 17292
rect 22189 17283 22247 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 25130 17280 25136 17332
rect 25188 17280 25194 17332
rect 25409 17323 25467 17329
rect 25409 17289 25421 17323
rect 25455 17320 25467 17323
rect 25590 17320 25596 17332
rect 25455 17292 25596 17320
rect 25455 17289 25467 17292
rect 25409 17283 25467 17289
rect 25590 17280 25596 17292
rect 25648 17280 25654 17332
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 19760 17224 20453 17252
rect 19760 17212 19766 17224
rect 20441 17221 20453 17224
rect 20487 17221 20499 17255
rect 20441 17215 20499 17221
rect 20533 17255 20591 17261
rect 20533 17221 20545 17255
rect 20579 17252 20591 17255
rect 20579 17224 21404 17252
rect 20579 17221 20591 17224
rect 20533 17215 20591 17221
rect 20254 17144 20260 17196
rect 20312 17144 20318 17196
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 20898 17184 20904 17196
rect 20772 17156 20904 17184
rect 20772 17144 20778 17156
rect 20898 17144 20904 17156
rect 20956 17184 20962 17196
rect 21177 17187 21235 17193
rect 21177 17184 21189 17187
rect 20956 17156 21189 17184
rect 20956 17144 20962 17156
rect 21177 17153 21189 17156
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 21266 17144 21272 17196
rect 21324 17184 21330 17196
rect 21376 17184 21404 17224
rect 22278 17212 22284 17264
rect 22336 17212 22342 17264
rect 21324 17156 21404 17184
rect 21324 17144 21330 17156
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21692 17156 21833 17184
rect 21692 17144 21698 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22002 17144 22008 17196
rect 22060 17144 22066 17196
rect 23290 17144 23296 17196
rect 23348 17144 23354 17196
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17153 23535 17187
rect 23477 17147 23535 17153
rect 19291 17088 19656 17116
rect 20073 17119 20131 17125
rect 19291 17085 19303 17088
rect 19245 17079 19303 17085
rect 20073 17085 20085 17119
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 17865 17051 17923 17057
rect 17865 17048 17877 17051
rect 15948 17020 17877 17048
rect 15565 17011 15623 17017
rect 17865 17017 17877 17020
rect 17911 17017 17923 17051
rect 17865 17011 17923 17017
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 20088 17048 20116 17079
rect 21082 17076 21088 17128
rect 21140 17076 21146 17128
rect 21358 17076 21364 17128
rect 21416 17076 21422 17128
rect 23014 17076 23020 17128
rect 23072 17076 23078 17128
rect 18564 17020 20116 17048
rect 18564 17008 18570 17020
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 22186 17048 22192 17060
rect 20588 17020 22192 17048
rect 20588 17008 20594 17020
rect 22186 17008 22192 17020
rect 22244 17048 22250 17060
rect 23492 17048 23520 17147
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 24026 17193 24032 17196
rect 24020 17184 24032 17193
rect 23987 17156 24032 17184
rect 24020 17147 24032 17156
rect 24026 17144 24032 17147
rect 24084 17144 24090 17196
rect 25148 17184 25176 17280
rect 25225 17187 25283 17193
rect 25225 17184 25237 17187
rect 25148 17156 25237 17184
rect 25225 17153 25237 17156
rect 25271 17153 25283 17187
rect 25225 17147 25283 17153
rect 25593 17187 25651 17193
rect 25593 17153 25605 17187
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25608 17116 25636 17147
rect 24820 17088 25636 17116
rect 24820 17076 24826 17088
rect 22244 17020 23520 17048
rect 22244 17008 22250 17020
rect 25774 17008 25780 17060
rect 25832 17008 25838 17060
rect 12308 16952 12756 16980
rect 12308 16940 12314 16952
rect 12894 16940 12900 16992
rect 12952 16940 12958 16992
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16980 14151 16983
rect 14550 16980 14556 16992
rect 14139 16952 14556 16980
rect 14139 16949 14151 16952
rect 14093 16943 14151 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 18690 16940 18696 16992
rect 18748 16940 18754 16992
rect 20806 16940 20812 16992
rect 20864 16940 20870 16992
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21876 16952 22017 16980
rect 21876 16940 21882 16952
rect 22005 16949 22017 16952
rect 22051 16980 22063 16983
rect 22462 16980 22468 16992
rect 22051 16952 22468 16980
rect 22051 16949 22063 16952
rect 22005 16943 22063 16949
rect 22462 16940 22468 16952
rect 22520 16980 22526 16992
rect 23290 16980 23296 16992
rect 22520 16952 23296 16980
rect 22520 16940 22526 16952
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 23661 16983 23719 16989
rect 23661 16980 23673 16983
rect 23624 16952 23673 16980
rect 23624 16940 23630 16952
rect 23661 16949 23673 16952
rect 23707 16949 23719 16983
rect 23661 16943 23719 16949
rect 1104 16890 26220 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 26220 16890
rect 1104 16816 26220 16838
rect 11790 16736 11796 16788
rect 11848 16736 11854 16788
rect 15930 16736 15936 16788
rect 15988 16776 15994 16788
rect 16209 16779 16267 16785
rect 16209 16776 16221 16779
rect 15988 16748 16221 16776
rect 15988 16736 15994 16748
rect 16209 16745 16221 16748
rect 16255 16745 16267 16779
rect 16209 16739 16267 16745
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 18506 16776 18512 16788
rect 18371 16748 18512 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16776 19947 16779
rect 20254 16776 20260 16788
rect 19935 16748 20260 16776
rect 19935 16745 19947 16748
rect 19889 16739 19947 16745
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 5626 16668 5632 16720
rect 5684 16708 5690 16720
rect 6638 16708 6644 16720
rect 5684 16680 6644 16708
rect 5684 16668 5690 16680
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 22152 16680 23612 16708
rect 22152 16668 22158 16680
rect 12250 16600 12256 16652
rect 12308 16600 12314 16652
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 6178 16532 6184 16584
rect 6236 16532 6242 16584
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 12360 16572 12388 16603
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12492 16612 13461 16640
rect 12492 16600 12498 16612
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13630 16600 13636 16652
rect 13688 16640 13694 16652
rect 15194 16640 15200 16652
rect 13688 16612 15200 16640
rect 13688 16600 13694 16612
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15344 16612 15577 16640
rect 15344 16600 15350 16612
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 16850 16640 16856 16652
rect 15795 16612 16856 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 16942 16600 16948 16652
rect 17000 16600 17006 16652
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 18380 16612 19257 16640
rect 18380 16600 18386 16612
rect 19245 16609 19257 16612
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20898 16640 20904 16652
rect 20303 16612 20904 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 23584 16649 23612 16680
rect 23569 16643 23627 16649
rect 21652 16612 21956 16640
rect 13648 16572 13676 16600
rect 12360 16544 13676 16572
rect 17212 16575 17270 16581
rect 17212 16541 17224 16575
rect 17258 16572 17270 16575
rect 18690 16572 18696 16584
rect 17258 16544 18696 16572
rect 17258 16541 17270 16544
rect 17212 16535 17270 16541
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19978 16532 19984 16584
rect 20036 16532 20042 16584
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20346 16572 20352 16584
rect 20119 16544 20352 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20346 16532 20352 16544
rect 20404 16532 20410 16584
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16572 21511 16575
rect 21652 16572 21680 16612
rect 21499 16544 21680 16572
rect 21729 16575 21787 16581
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 12161 16507 12219 16513
rect 12161 16473 12173 16507
rect 12207 16504 12219 16507
rect 12207 16476 12434 16504
rect 12207 16473 12219 16476
rect 12161 16467 12219 16473
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 11606 16436 11612 16448
rect 1636 16408 11612 16436
rect 1636 16396 1642 16408
rect 11606 16396 11612 16408
rect 11664 16396 11670 16448
rect 12406 16436 12434 16476
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 19150 16504 19156 16516
rect 13044 16476 19156 16504
rect 13044 16464 13050 16476
rect 19150 16464 19156 16476
rect 19208 16464 19214 16516
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 20257 16507 20315 16513
rect 20257 16504 20269 16507
rect 19760 16476 20269 16504
rect 19760 16464 19766 16476
rect 20257 16473 20269 16476
rect 20303 16473 20315 16507
rect 20824 16504 20852 16535
rect 20898 16504 20904 16516
rect 20824 16476 20904 16504
rect 20257 16467 20315 16473
rect 20898 16464 20904 16476
rect 20956 16464 20962 16516
rect 21266 16464 21272 16516
rect 21324 16504 21330 16516
rect 21744 16504 21772 16535
rect 21818 16532 21824 16584
rect 21876 16532 21882 16584
rect 21928 16572 21956 16612
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 22097 16575 22155 16581
rect 22097 16572 22109 16575
rect 21928 16544 22109 16572
rect 22097 16541 22109 16544
rect 22143 16541 22155 16575
rect 23014 16572 23020 16584
rect 22097 16535 22155 16541
rect 22296 16544 23020 16572
rect 21324 16476 21772 16504
rect 21324 16464 21330 16476
rect 21910 16464 21916 16516
rect 21968 16464 21974 16516
rect 22296 16513 22324 16544
rect 23014 16532 23020 16544
rect 23072 16572 23078 16584
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 23072 16544 24409 16572
rect 23072 16532 23078 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 22281 16507 22339 16513
rect 22281 16473 22293 16507
rect 22327 16473 22339 16507
rect 24642 16507 24700 16513
rect 24642 16504 24654 16507
rect 22281 16467 22339 16473
rect 24228 16476 24654 16504
rect 12802 16436 12808 16448
rect 12406 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 12894 16396 12900 16448
rect 12952 16396 12958 16448
rect 15838 16396 15844 16448
rect 15896 16396 15902 16448
rect 20533 16439 20591 16445
rect 20533 16405 20545 16439
rect 20579 16436 20591 16439
rect 21082 16436 21088 16448
rect 20579 16408 21088 16436
rect 20579 16405 20591 16408
rect 20533 16399 20591 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 21542 16396 21548 16448
rect 21600 16396 21606 16448
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 22296 16436 22324 16467
rect 21784 16408 22324 16436
rect 21784 16396 21790 16408
rect 23750 16396 23756 16448
rect 23808 16396 23814 16448
rect 23842 16396 23848 16448
rect 23900 16396 23906 16448
rect 24228 16445 24256 16476
rect 24642 16473 24654 16476
rect 24688 16473 24700 16507
rect 24642 16467 24700 16473
rect 24213 16439 24271 16445
rect 24213 16405 24225 16439
rect 24259 16405 24271 16439
rect 24213 16399 24271 16405
rect 25498 16396 25504 16448
rect 25556 16436 25562 16448
rect 25777 16439 25835 16445
rect 25777 16436 25789 16439
rect 25556 16408 25789 16436
rect 25556 16396 25562 16408
rect 25777 16405 25789 16408
rect 25823 16405 25835 16439
rect 25777 16399 25835 16405
rect 1104 16346 26220 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 26220 16346
rect 1104 16272 26220 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 4433 16235 4491 16241
rect 4433 16201 4445 16235
rect 4479 16232 4491 16235
rect 4614 16232 4620 16244
rect 4479 16204 4620 16232
rect 4479 16201 4491 16204
rect 4433 16195 4491 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 5868 16204 6101 16232
rect 5868 16192 5874 16204
rect 6089 16201 6101 16204
rect 6135 16201 6147 16235
rect 6089 16195 6147 16201
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 12492 16204 12909 16232
rect 12492 16192 12498 16204
rect 12897 16201 12909 16204
rect 12943 16201 12955 16235
rect 12897 16195 12955 16201
rect 18322 16192 18328 16244
rect 18380 16192 18386 16244
rect 20806 16232 20812 16244
rect 18984 16204 20812 16232
rect 1762 16124 1768 16176
rect 1820 16164 1826 16176
rect 1820 16136 5488 16164
rect 1820 16124 1826 16136
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 2314 16056 2320 16108
rect 2372 16056 2378 16108
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 2573 16099 2631 16105
rect 2573 16096 2585 16099
rect 2464 16068 2585 16096
rect 2464 16056 2470 16068
rect 2573 16065 2585 16068
rect 2619 16065 2631 16099
rect 2573 16059 2631 16065
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3936 16068 3985 16096
rect 3936 16056 3942 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4492 16099 4550 16105
rect 4492 16065 4504 16099
rect 4538 16096 4550 16099
rect 4798 16096 4804 16108
rect 4538 16068 4804 16096
rect 4538 16065 4550 16068
rect 4492 16059 4550 16065
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 3697 15895 3755 15901
rect 3697 15861 3709 15895
rect 3743 15892 3755 15895
rect 4062 15892 4068 15904
rect 3743 15864 4068 15892
rect 3743 15861 3755 15864
rect 3697 15855 3755 15861
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4706 15892 4712 15904
rect 4663 15864 4712 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 5460 15892 5488 16136
rect 5534 16124 5540 16176
rect 5592 16164 5598 16176
rect 5629 16167 5687 16173
rect 5629 16164 5641 16167
rect 5592 16136 5641 16164
rect 5592 16124 5598 16136
rect 5629 16133 5641 16136
rect 5675 16164 5687 16167
rect 6178 16164 6184 16176
rect 5675 16136 6184 16164
rect 5675 16133 5687 16136
rect 5629 16127 5687 16133
rect 6178 16124 6184 16136
rect 6236 16164 6242 16176
rect 6549 16167 6607 16173
rect 6549 16164 6561 16167
rect 6236 16136 6561 16164
rect 6236 16124 6242 16136
rect 6549 16133 6561 16136
rect 6595 16133 6607 16167
rect 6549 16127 6607 16133
rect 11698 16124 11704 16176
rect 11756 16164 11762 16176
rect 17212 16167 17270 16173
rect 11756 16136 14412 16164
rect 11756 16124 11762 16136
rect 6362 16096 6368 16108
rect 5920 16068 6368 16096
rect 5920 15972 5948 16068
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 11784 16099 11842 16105
rect 11784 16065 11796 16099
rect 11830 16096 11842 16099
rect 12066 16096 12072 16108
rect 11830 16068 12072 16096
rect 11830 16065 11842 16068
rect 11784 16059 11842 16065
rect 12066 16056 12072 16068
rect 12124 16056 12130 16108
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 14384 16105 14412 16136
rect 17212 16133 17224 16167
rect 17258 16164 17270 16167
rect 18984 16164 19012 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 22833 16235 22891 16241
rect 22833 16201 22845 16235
rect 22879 16232 22891 16235
rect 23750 16232 23756 16244
rect 22879 16204 23756 16232
rect 22879 16201 22891 16204
rect 22833 16195 22891 16201
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 23842 16192 23848 16244
rect 23900 16232 23906 16244
rect 24857 16235 24915 16241
rect 24857 16232 24869 16235
rect 23900 16204 24869 16232
rect 23900 16192 23906 16204
rect 24857 16201 24869 16204
rect 24903 16201 24915 16235
rect 24857 16195 24915 16201
rect 22465 16167 22523 16173
rect 17258 16136 19012 16164
rect 19996 16136 21680 16164
rect 17258 16133 17270 16136
rect 17212 16127 17270 16133
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 13495 16068 13829 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 14369 16099 14427 16105
rect 14369 16065 14381 16099
rect 14415 16065 14427 16099
rect 14369 16059 14427 16065
rect 16942 16056 16948 16108
rect 17000 16056 17006 16108
rect 19702 16056 19708 16108
rect 19760 16105 19766 16108
rect 19996 16105 20024 16136
rect 19760 16096 19772 16105
rect 19981 16099 20039 16105
rect 19760 16068 19805 16096
rect 19760 16059 19772 16068
rect 19981 16065 19993 16099
rect 20027 16065 20039 16099
rect 20898 16096 20904 16108
rect 19981 16059 20039 16065
rect 20272 16068 20904 16096
rect 19760 16056 19766 16059
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11020 16000 11529 16028
rect 11020 15988 11026 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 13630 15988 13636 16040
rect 13688 15988 13694 16040
rect 5902 15920 5908 15972
rect 5960 15920 5966 15972
rect 12989 15963 13047 15969
rect 12989 15960 13001 15963
rect 6472 15932 11560 15960
rect 6472 15892 6500 15932
rect 5460 15864 6500 15892
rect 6546 15852 6552 15904
rect 6604 15892 6610 15904
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 6604 15864 6745 15892
rect 6604 15852 6610 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 11532 15892 11560 15932
rect 12728 15932 13001 15960
rect 11790 15892 11796 15904
rect 11532 15864 11796 15892
rect 6733 15855 6791 15861
rect 11790 15852 11796 15864
rect 11848 15852 11854 15904
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12728 15892 12756 15932
rect 12989 15929 13001 15932
rect 13035 15929 13047 15963
rect 12989 15923 13047 15929
rect 20272 15904 20300 16068
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 21381 16099 21439 16105
rect 21381 16065 21393 16099
rect 21427 16096 21439 16099
rect 21542 16096 21548 16108
rect 21427 16068 21548 16096
rect 21427 16065 21439 16068
rect 21381 16059 21439 16065
rect 21542 16056 21548 16068
rect 21600 16056 21606 16108
rect 21652 16037 21680 16136
rect 22465 16133 22477 16167
rect 22511 16164 22523 16167
rect 23014 16164 23020 16176
rect 22511 16136 23020 16164
rect 22511 16133 22523 16136
rect 22465 16127 22523 16133
rect 23014 16124 23020 16136
rect 23072 16164 23078 16176
rect 23109 16167 23167 16173
rect 23109 16164 23121 16167
rect 23072 16136 23121 16164
rect 23072 16124 23078 16136
rect 23109 16133 23121 16136
rect 23155 16164 23167 16167
rect 23155 16136 23796 16164
rect 23155 16133 23167 16136
rect 23109 16127 23167 16133
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16065 21879 16099
rect 21821 16059 21879 16065
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 16028 21695 16031
rect 21726 16028 21732 16040
rect 21683 16000 21732 16028
rect 21683 15997 21695 16000
rect 21637 15991 21695 15997
rect 21726 15988 21732 16000
rect 21784 15988 21790 16040
rect 12308 15864 12756 15892
rect 12308 15852 12314 15864
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 17862 15892 17868 15904
rect 15344 15864 17868 15892
rect 15344 15852 15350 15864
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 18601 15895 18659 15901
rect 18601 15861 18613 15895
rect 18647 15892 18659 15895
rect 18690 15892 18696 15904
rect 18647 15864 18696 15892
rect 18647 15861 18659 15864
rect 18601 15855 18659 15861
rect 18690 15852 18696 15864
rect 18748 15852 18754 15904
rect 20254 15852 20260 15904
rect 20312 15852 20318 15904
rect 20346 15852 20352 15904
rect 20404 15892 20410 15904
rect 21836 15892 21864 16059
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22281 16099 22339 16105
rect 22281 16096 22293 16099
rect 22152 16068 22293 16096
rect 22152 16056 22158 16068
rect 22281 16065 22293 16068
rect 22327 16065 22339 16099
rect 22281 16059 22339 16065
rect 22554 16056 22560 16108
rect 22612 16056 22618 16108
rect 22646 16056 22652 16108
rect 22704 16056 22710 16108
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16065 22983 16099
rect 22925 16059 22983 16065
rect 21913 16031 21971 16037
rect 21913 15997 21925 16031
rect 21959 16028 21971 16031
rect 22940 16028 22968 16059
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 23308 16028 23336 16059
rect 23566 16056 23572 16108
rect 23624 16056 23630 16108
rect 23768 16105 23796 16136
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 23842 16056 23848 16108
rect 23900 16056 23906 16108
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16065 23995 16099
rect 23937 16059 23995 16065
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 25498 16096 25504 16108
rect 24627 16068 25504 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 23952 16028 23980 16059
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16096 25651 16099
rect 25682 16096 25688 16108
rect 25639 16068 25688 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 21959 16000 22968 16028
rect 23216 16000 23980 16028
rect 21959 15997 21971 16000
rect 21913 15991 21971 15997
rect 22646 15920 22652 15972
rect 22704 15960 22710 15972
rect 23106 15960 23112 15972
rect 22704 15932 23112 15960
rect 22704 15920 22710 15932
rect 23106 15920 23112 15932
rect 23164 15960 23170 15972
rect 23216 15960 23244 16000
rect 23164 15932 23244 15960
rect 24121 15963 24179 15969
rect 23164 15920 23170 15932
rect 24121 15929 24133 15963
rect 24167 15960 24179 15963
rect 24486 15960 24492 15972
rect 24167 15932 24492 15960
rect 24167 15929 24179 15932
rect 24121 15923 24179 15929
rect 24486 15920 24492 15932
rect 24544 15920 24550 15972
rect 24762 15920 24768 15972
rect 24820 15920 24826 15972
rect 20404 15864 21864 15892
rect 23477 15895 23535 15901
rect 20404 15852 20410 15864
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 24578 15892 24584 15904
rect 23523 15864 24584 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 25774 15852 25780 15904
rect 25832 15852 25838 15904
rect 1104 15802 26220 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 26220 15802
rect 1104 15728 26220 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 1762 15688 1768 15700
rect 1627 15660 1768 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 2406 15648 2412 15700
rect 2464 15648 2470 15700
rect 2590 15648 2596 15700
rect 2648 15648 2654 15700
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6788 15660 6929 15688
rect 6788 15648 6794 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 10965 15691 11023 15697
rect 10965 15657 10977 15691
rect 11011 15688 11023 15691
rect 11698 15688 11704 15700
rect 11011 15660 11704 15688
rect 11011 15657 11023 15660
rect 10965 15651 11023 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 12124 15660 12449 15688
rect 12124 15648 12130 15660
rect 12437 15657 12449 15660
rect 12483 15657 12495 15691
rect 12437 15651 12495 15657
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 18233 15691 18291 15697
rect 18233 15688 18245 15691
rect 13412 15660 18245 15688
rect 13412 15648 13418 15660
rect 18233 15657 18245 15660
rect 18279 15657 18291 15691
rect 18233 15651 18291 15657
rect 20165 15691 20223 15697
rect 20165 15657 20177 15691
rect 20211 15688 20223 15691
rect 21358 15688 21364 15700
rect 20211 15660 21364 15688
rect 20211 15657 20223 15660
rect 20165 15651 20223 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 22281 15691 22339 15697
rect 22281 15657 22293 15691
rect 22327 15688 22339 15691
rect 23750 15688 23756 15700
rect 22327 15660 23756 15688
rect 22327 15657 22339 15660
rect 22281 15651 22339 15657
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 25777 15691 25835 15697
rect 25777 15657 25789 15691
rect 25823 15688 25835 15691
rect 26050 15688 26056 15700
rect 25823 15660 26056 15688
rect 25823 15657 25835 15660
rect 25777 15651 25835 15657
rect 26050 15648 26056 15660
rect 26108 15648 26114 15700
rect 12802 15580 12808 15632
rect 12860 15620 12866 15632
rect 17405 15623 17463 15629
rect 17405 15620 17417 15623
rect 12860 15592 17417 15620
rect 12860 15580 12866 15592
rect 17405 15589 17417 15592
rect 17451 15589 17463 15623
rect 18506 15620 18512 15632
rect 17405 15583 17463 15589
rect 17880 15592 18512 15620
rect 3234 15552 3240 15564
rect 2746 15524 3240 15552
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 2746 15484 2774 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3326 15512 3332 15564
rect 3384 15552 3390 15564
rect 5902 15552 5908 15564
rect 3384 15524 4384 15552
rect 3384 15512 3390 15524
rect 2363 15456 2774 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 1486 15376 1492 15428
rect 1544 15376 1550 15428
rect 2148 15348 2176 15447
rect 2866 15444 2872 15496
rect 2924 15444 2930 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3602 15484 3608 15496
rect 3099 15456 3608 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 4062 15444 4068 15496
rect 4120 15444 4126 15496
rect 2225 15419 2283 15425
rect 2225 15385 2237 15419
rect 2271 15416 2283 15419
rect 2561 15419 2619 15425
rect 2561 15416 2573 15419
rect 2271 15388 2573 15416
rect 2271 15385 2283 15388
rect 2225 15379 2283 15385
rect 2561 15385 2573 15388
rect 2607 15385 2619 15419
rect 2561 15379 2619 15385
rect 2682 15376 2688 15428
rect 2740 15416 2746 15428
rect 2777 15419 2835 15425
rect 2777 15416 2789 15419
rect 2740 15388 2789 15416
rect 2740 15376 2746 15388
rect 2777 15385 2789 15388
rect 2823 15385 2835 15419
rect 2777 15379 2835 15385
rect 3326 15376 3332 15428
rect 3384 15376 3390 15428
rect 3513 15419 3571 15425
rect 3513 15385 3525 15419
rect 3559 15416 3571 15419
rect 3970 15416 3976 15428
rect 3559 15388 3976 15416
rect 3559 15385 3571 15388
rect 3513 15379 3571 15385
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 4356 15425 4384 15524
rect 5643 15524 5908 15552
rect 5643 15493 5671 15524
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 9508 15524 10272 15552
rect 5628 15487 5686 15493
rect 5628 15453 5640 15487
rect 5674 15453 5686 15487
rect 5628 15447 5686 15453
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15484 6791 15487
rect 7374 15484 7380 15496
rect 6779 15456 7380 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 4341 15419 4399 15425
rect 4341 15385 4353 15419
rect 4387 15416 4399 15419
rect 5736 15416 5764 15444
rect 4387 15388 5764 15416
rect 4387 15385 4399 15388
rect 4341 15379 4399 15385
rect 6748 15360 6776 15447
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 8570 15444 8576 15496
rect 8628 15484 8634 15496
rect 9508 15493 9536 15524
rect 10244 15493 10272 15524
rect 12894 15512 12900 15564
rect 12952 15512 12958 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13630 15552 13636 15564
rect 13127 15524 13636 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 15013 15555 15071 15561
rect 15013 15552 15025 15555
rect 14844 15524 15025 15552
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 8628 15456 9505 15484
rect 8628 15444 8634 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9493 15447 9551 15453
rect 9876 15456 10057 15484
rect 9030 15376 9036 15428
rect 9088 15416 9094 15428
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 9088 15388 9321 15416
rect 9088 15376 9094 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9309 15379 9367 15385
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 9876 15425 9904 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 12089 15487 12147 15493
rect 12089 15453 12101 15487
rect 12135 15484 12147 15487
rect 12250 15484 12256 15496
rect 12135 15456 12256 15484
rect 12135 15453 12147 15456
rect 12089 15447 12147 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 14844 15484 14872 15524
rect 15013 15521 15025 15524
rect 15059 15552 15071 15555
rect 15286 15552 15292 15564
rect 15059 15524 15292 15552
rect 15059 15521 15071 15524
rect 15013 15515 15071 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15378 15512 15384 15564
rect 15436 15512 15442 15564
rect 17880 15561 17908 15592
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 20346 15580 20352 15632
rect 20404 15620 20410 15632
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20404 15592 20637 15620
rect 20404 15580 20410 15592
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 22465 15623 22523 15629
rect 22465 15620 22477 15623
rect 20625 15583 20683 15589
rect 21652 15592 22477 15620
rect 17865 15555 17923 15561
rect 17865 15521 17877 15555
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 21652 15561 21680 15592
rect 22465 15589 22477 15592
rect 22511 15620 22523 15623
rect 22646 15620 22652 15632
rect 22511 15592 22652 15620
rect 22511 15589 22523 15592
rect 22465 15583 22523 15589
rect 22646 15580 22652 15592
rect 22704 15580 22710 15632
rect 24213 15623 24271 15629
rect 24213 15589 24225 15623
rect 24259 15620 24271 15623
rect 24259 15592 24992 15620
rect 24259 15589 24271 15592
rect 24213 15583 24271 15589
rect 24964 15564 24992 15592
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18012 15524 18797 15552
rect 18012 15512 18018 15524
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 21637 15555 21695 15561
rect 21637 15521 21649 15555
rect 21683 15521 21695 15555
rect 21637 15515 21695 15521
rect 21726 15512 21732 15564
rect 21784 15552 21790 15564
rect 22738 15552 22744 15564
rect 21784 15524 22744 15552
rect 21784 15512 21790 15524
rect 22738 15512 22744 15524
rect 22796 15552 22802 15564
rect 22833 15555 22891 15561
rect 22833 15552 22845 15555
rect 22796 15524 22845 15552
rect 22796 15512 22802 15524
rect 22833 15521 22845 15524
rect 22879 15521 22891 15555
rect 22833 15515 22891 15521
rect 24946 15512 24952 15564
rect 25004 15512 25010 15564
rect 13228 15456 14872 15484
rect 14921 15487 14979 15493
rect 13228 15444 13234 15456
rect 14921 15453 14933 15487
rect 14967 15484 14979 15487
rect 14967 15456 18644 15484
rect 14967 15453 14979 15456
rect 14921 15447 14979 15453
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 9640 15388 9873 15416
rect 9640 15376 9646 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9861 15379 9919 15385
rect 12805 15419 12863 15425
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 12851 15388 13584 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 2958 15348 2964 15360
rect 2148 15320 2964 15348
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3142 15308 3148 15360
rect 3200 15308 3206 15360
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 4798 15348 4804 15360
rect 4203 15320 4804 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 5350 15308 5356 15360
rect 5408 15308 5414 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 6730 15348 6736 15360
rect 6503 15320 6736 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9769 15351 9827 15357
rect 9769 15348 9781 15351
rect 8996 15320 9781 15348
rect 8996 15308 9002 15320
rect 9769 15317 9781 15320
rect 9815 15317 9827 15351
rect 9769 15311 9827 15317
rect 10226 15308 10232 15360
rect 10284 15308 10290 15360
rect 13354 15308 13360 15360
rect 13412 15308 13418 15360
rect 13556 15348 13584 15388
rect 13630 15376 13636 15428
rect 13688 15376 13694 15428
rect 17773 15419 17831 15425
rect 17773 15385 17785 15419
rect 17819 15416 17831 15419
rect 18506 15416 18512 15428
rect 17819 15388 18512 15416
rect 17819 15385 17831 15388
rect 17773 15379 17831 15385
rect 18506 15376 18512 15388
rect 18564 15376 18570 15428
rect 18616 15416 18644 15456
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 18748 15456 19349 15484
rect 18748 15444 18754 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 19981 15487 20039 15493
rect 19981 15453 19993 15487
rect 20027 15484 20039 15487
rect 20073 15487 20131 15493
rect 20073 15484 20085 15487
rect 20027 15456 20085 15484
rect 20027 15453 20039 15456
rect 19981 15447 20039 15453
rect 20073 15453 20085 15456
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20220 15456 20545 15484
rect 20220 15444 20226 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20714 15444 20720 15496
rect 20772 15444 20778 15496
rect 21910 15444 21916 15496
rect 21968 15444 21974 15496
rect 22646 15444 22652 15496
rect 22704 15484 22710 15496
rect 23658 15484 23664 15496
rect 22704 15456 23664 15484
rect 22704 15444 22710 15456
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 25222 15444 25228 15496
rect 25280 15444 25286 15496
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15453 25651 15487
rect 25593 15447 25651 15453
rect 20254 15416 20260 15428
rect 18616 15388 20260 15416
rect 20254 15376 20260 15388
rect 20312 15376 20318 15428
rect 23100 15419 23158 15425
rect 23100 15385 23112 15419
rect 23146 15416 23158 15419
rect 23290 15416 23296 15428
rect 23146 15388 23296 15416
rect 23146 15385 23158 15388
rect 23100 15379 23158 15385
rect 23290 15376 23296 15388
rect 23348 15376 23354 15428
rect 23382 15376 23388 15428
rect 23440 15416 23446 15428
rect 25608 15416 25636 15447
rect 23440 15388 25636 15416
rect 23440 15376 23446 15388
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 13556 15320 14473 15348
rect 14461 15317 14473 15320
rect 14507 15317 14519 15351
rect 14461 15311 14519 15317
rect 14826 15308 14832 15360
rect 14884 15308 14890 15360
rect 15930 15308 15936 15360
rect 15988 15308 15994 15360
rect 18598 15308 18604 15360
rect 18656 15308 18662 15360
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 21821 15351 21879 15357
rect 21821 15348 21833 15351
rect 21048 15320 21833 15348
rect 21048 15308 21054 15320
rect 21821 15317 21833 15320
rect 21867 15317 21879 15351
rect 21821 15311 21879 15317
rect 24302 15308 24308 15360
rect 24360 15348 24366 15360
rect 24397 15351 24455 15357
rect 24397 15348 24409 15351
rect 24360 15320 24409 15348
rect 24360 15308 24366 15320
rect 24397 15317 24409 15320
rect 24443 15317 24455 15351
rect 24397 15311 24455 15317
rect 25406 15308 25412 15360
rect 25464 15308 25470 15360
rect 1104 15258 26220 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 26220 15258
rect 1104 15184 26220 15206
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 3142 15144 3148 15156
rect 2823 15116 3148 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 4433 15147 4491 15153
rect 4433 15144 4445 15147
rect 4028 15116 4445 15144
rect 4028 15104 4034 15116
rect 4433 15113 4445 15116
rect 4479 15113 4491 15147
rect 5534 15144 5540 15156
rect 4433 15107 4491 15113
rect 5000 15116 5540 15144
rect 1949 15079 2007 15085
rect 1949 15045 1961 15079
rect 1995 15045 2007 15079
rect 1949 15039 2007 15045
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15076 3019 15079
rect 3298 15079 3356 15085
rect 3298 15076 3310 15079
rect 3007 15048 3310 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 3298 15045 3310 15048
rect 3344 15045 3356 15079
rect 4448 15076 4476 15107
rect 4448 15048 4660 15076
rect 3298 15039 3356 15045
rect 1964 15008 1992 15039
rect 2590 15008 2596 15020
rect 1964 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 2866 15008 2872 15020
rect 2731 14980 2872 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 2866 14968 2872 14980
rect 2924 15008 2930 15020
rect 3142 15008 3148 15020
rect 2924 14980 3148 15008
rect 2924 14968 2930 14980
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4212 14980 4537 15008
rect 4212 14968 4218 14980
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 1964 14912 2452 14940
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14804 1823 14807
rect 1854 14804 1860 14816
rect 1811 14776 1860 14804
rect 1811 14773 1823 14776
rect 1765 14767 1823 14773
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 1964 14813 1992 14912
rect 2424 14881 2452 14912
rect 3050 14900 3056 14952
rect 3108 14900 3114 14952
rect 4632 14940 4660 15048
rect 5000 15017 5028 15116
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 13262 15144 13268 15156
rect 12299 15116 13268 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 15565 15147 15623 15153
rect 13412 15116 15516 15144
rect 13412 15104 13418 15116
rect 5077 15079 5135 15085
rect 5077 15045 5089 15079
rect 5123 15076 5135 15079
rect 5123 15048 5304 15076
rect 5123 15045 5135 15048
rect 5077 15039 5135 15045
rect 5276 15017 5304 15048
rect 5350 15036 5356 15088
rect 5408 15076 5414 15088
rect 5445 15079 5503 15085
rect 5445 15076 5457 15079
rect 5408 15048 5457 15076
rect 5408 15036 5414 15048
rect 5445 15045 5457 15048
rect 5491 15045 5503 15079
rect 5445 15039 5503 15045
rect 5810 15036 5816 15088
rect 5868 15076 5874 15088
rect 6365 15079 6423 15085
rect 6365 15076 6377 15079
rect 5868 15048 6377 15076
rect 5868 15036 5874 15048
rect 6365 15045 6377 15048
rect 6411 15045 6423 15079
rect 10962 15076 10968 15088
rect 6365 15039 6423 15045
rect 9968 15048 10968 15076
rect 4985 15011 5043 15017
rect 4985 14977 4997 15011
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 5994 15008 6000 15020
rect 5675 14980 6000 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5184 14940 5212 14971
rect 5552 14940 5580 14971
rect 5994 14968 6000 14980
rect 6052 15008 6058 15020
rect 6638 15008 6644 15020
rect 6052 14980 6644 15008
rect 6052 14968 6058 14980
rect 6638 14968 6644 14980
rect 6696 14968 6702 15020
rect 6733 15011 6791 15017
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7650 15008 7656 15020
rect 6779 14980 7656 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 7650 14968 7656 14980
rect 7708 15008 7714 15020
rect 9122 15008 9128 15020
rect 7708 14980 9128 15008
rect 7708 14968 7714 14980
rect 4632 14912 5580 14940
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 6549 14943 6607 14949
rect 6549 14940 6561 14943
rect 5776 14912 6561 14940
rect 5776 14900 5782 14912
rect 6549 14909 6561 14912
rect 6595 14909 6607 14943
rect 6549 14903 6607 14909
rect 2317 14875 2375 14881
rect 2317 14841 2329 14875
rect 2363 14841 2375 14875
rect 2317 14835 2375 14841
rect 2409 14875 2467 14881
rect 2409 14841 2421 14875
rect 2455 14872 2467 14875
rect 2682 14872 2688 14884
rect 2455 14844 2688 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 1949 14807 2007 14813
rect 1949 14773 1961 14807
rect 1995 14773 2007 14807
rect 2332 14804 2360 14835
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 6638 14832 6644 14884
rect 6696 14832 6702 14884
rect 8496 14881 8524 14980
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9594 15011 9652 15017
rect 9594 15008 9606 15011
rect 9272 14980 9606 15008
rect 9272 14968 9278 14980
rect 9594 14977 9606 14980
rect 9640 14977 9652 15011
rect 9594 14971 9652 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9968 15017 9996 15048
rect 10962 15036 10968 15048
rect 11020 15076 11026 15088
rect 12342 15076 12348 15088
rect 11020 15048 12348 15076
rect 11020 15036 11026 15048
rect 12342 15036 12348 15048
rect 12400 15076 12406 15088
rect 12400 15048 13676 15076
rect 12400 15036 12406 15048
rect 10226 15017 10232 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9824 14980 9873 15008
rect 9824 14968 9830 14980
rect 9861 14977 9873 14980
rect 9907 15008 9919 15011
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9907 14980 9965 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 9953 14977 9965 14980
rect 9999 14977 10011 15011
rect 10220 15008 10232 15017
rect 10187 14980 10232 15008
rect 9953 14971 10011 14977
rect 10220 14971 10232 14980
rect 10226 14968 10232 14971
rect 10284 14968 10290 15020
rect 11606 14968 11612 15020
rect 11664 14968 11670 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 12161 15011 12219 15017
rect 12161 14977 12173 15011
rect 12207 15008 12219 15011
rect 13078 15008 13084 15020
rect 12207 14980 13084 15008
rect 12207 14977 12219 14980
rect 12161 14971 12219 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13354 14968 13360 15020
rect 13412 15017 13418 15020
rect 13648 15017 13676 15048
rect 13998 15017 14004 15020
rect 13412 15008 13424 15017
rect 13633 15011 13691 15017
rect 13412 14980 13457 15008
rect 13412 14971 13424 14980
rect 13633 14977 13645 15011
rect 13679 15008 13691 15011
rect 13725 15011 13783 15017
rect 13725 15008 13737 15011
rect 13679 14980 13737 15008
rect 13679 14977 13691 14980
rect 13633 14971 13691 14977
rect 13725 14977 13737 14980
rect 13771 14977 13783 15011
rect 13725 14971 13783 14977
rect 13992 14971 14004 15017
rect 13412 14968 13418 14971
rect 13998 14968 14004 14971
rect 14056 14968 14062 15020
rect 15194 14900 15200 14952
rect 15252 14900 15258 14952
rect 15488 14940 15516 15116
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 15930 15144 15936 15156
rect 15611 15116 15936 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 15930 15104 15936 15116
rect 15988 15104 15994 15156
rect 22002 15104 22008 15156
rect 22060 15144 22066 15156
rect 22060 15116 22232 15144
rect 22060 15104 22066 15116
rect 15657 15079 15715 15085
rect 15657 15045 15669 15079
rect 15703 15076 15715 15079
rect 15746 15076 15752 15088
rect 15703 15048 15752 15076
rect 15703 15045 15715 15048
rect 15657 15039 15715 15045
rect 15746 15036 15752 15048
rect 15804 15036 15810 15088
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 17184 15048 18092 15076
rect 17184 15036 17190 15048
rect 18064 15017 18092 15048
rect 22094 15036 22100 15088
rect 22152 15036 22158 15088
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 15008 17095 15011
rect 17497 15011 17555 15017
rect 17497 15008 17509 15011
rect 17083 14980 17509 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17497 14977 17509 14980
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 22204 15017 22232 15116
rect 23290 15104 23296 15156
rect 23348 15104 23354 15156
rect 23661 15147 23719 15153
rect 23661 15113 23673 15147
rect 23707 15144 23719 15147
rect 24302 15144 24308 15156
rect 23707 15116 24308 15144
rect 23707 15113 23719 15116
rect 23661 15107 23719 15113
rect 24302 15104 24308 15116
rect 24360 15104 24366 15156
rect 25133 15147 25191 15153
rect 25133 15113 25145 15147
rect 25179 15144 25191 15147
rect 25222 15144 25228 15156
rect 25179 15116 25228 15144
rect 25179 15113 25191 15116
rect 25133 15107 25191 15113
rect 25222 15104 25228 15116
rect 25280 15104 25286 15156
rect 23750 15036 23756 15088
rect 23808 15036 23814 15088
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21508 14980 22017 15008
rect 21508 14968 21514 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 24946 14968 24952 15020
rect 25004 14968 25010 15020
rect 15749 14943 15807 14949
rect 15749 14940 15761 14943
rect 15488 14912 15761 14940
rect 15749 14909 15761 14912
rect 15795 14909 15807 14943
rect 15749 14903 15807 14909
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14841 8539 14875
rect 15212 14872 15240 14900
rect 15562 14872 15568 14884
rect 15212 14844 15568 14872
rect 8481 14835 8539 14841
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 15764 14872 15792 14903
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 16816 14912 17141 14940
rect 16816 14900 16822 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14909 17279 14943
rect 17221 14903 17279 14909
rect 17236 14872 17264 14903
rect 20438 14900 20444 14952
rect 20496 14940 20502 14952
rect 23845 14943 23903 14949
rect 20496 14912 22968 14940
rect 20496 14900 20502 14912
rect 15764 14844 17264 14872
rect 17310 14832 17316 14884
rect 17368 14872 17374 14884
rect 22646 14872 22652 14884
rect 17368 14844 22652 14872
rect 17368 14832 17374 14844
rect 22646 14832 22652 14844
rect 22704 14832 22710 14884
rect 22940 14872 22968 14912
rect 23845 14909 23857 14943
rect 23891 14909 23903 14943
rect 23845 14903 23903 14909
rect 23860 14872 23888 14903
rect 22940 14844 23888 14872
rect 2866 14804 2872 14816
rect 2332 14776 2872 14804
rect 1949 14767 2007 14773
rect 2866 14764 2872 14776
rect 2924 14804 2930 14816
rect 3326 14804 3332 14816
rect 2924 14776 3332 14804
rect 2924 14764 2930 14776
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 3752 14776 4629 14804
rect 3752 14764 3758 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 5626 14804 5632 14816
rect 5040 14776 5632 14804
rect 5040 14764 5046 14776
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 5813 14807 5871 14813
rect 5813 14773 5825 14807
rect 5859 14804 5871 14807
rect 6086 14804 6092 14816
rect 5859 14776 6092 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 11330 14764 11336 14816
rect 11388 14764 11394 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14826 14804 14832 14816
rect 13964 14776 14832 14804
rect 13964 14764 13970 14776
rect 14826 14764 14832 14776
rect 14884 14804 14890 14816
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 14884 14776 15117 14804
rect 14884 14764 14890 14776
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15105 14767 15163 14773
rect 15197 14807 15255 14813
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15378 14804 15384 14816
rect 15243 14776 15384 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 16666 14764 16672 14816
rect 16724 14764 16730 14816
rect 21726 14764 21732 14816
rect 21784 14804 21790 14816
rect 24854 14804 24860 14816
rect 21784 14776 24860 14804
rect 21784 14764 21790 14776
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 1104 14714 26220 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 26220 14714
rect 1104 14640 26220 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 3160 14532 3188 14563
rect 3234 14560 3240 14612
rect 3292 14560 3298 14612
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3694 14600 3700 14612
rect 3476 14572 3700 14600
rect 3476 14560 3482 14572
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 4798 14600 4804 14612
rect 4479 14572 4804 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 3326 14532 3332 14544
rect 3160 14504 3332 14532
rect 3326 14492 3332 14504
rect 3384 14532 3390 14544
rect 4448 14532 4476 14563
rect 4798 14560 4804 14572
rect 4856 14600 4862 14612
rect 5074 14600 5080 14612
rect 4856 14572 5080 14600
rect 4856 14560 4862 14572
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5184 14572 5641 14600
rect 3384 14504 4476 14532
rect 4617 14535 4675 14541
rect 3384 14492 3390 14504
rect 4617 14501 4629 14535
rect 4663 14501 4675 14535
rect 4617 14495 4675 14501
rect 3142 14424 3148 14476
rect 3200 14464 3206 14476
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3200 14436 3893 14464
rect 3200 14424 3206 14436
rect 1578 14356 1584 14408
rect 1636 14396 1642 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1636 14368 1777 14396
rect 1636 14356 1642 14368
rect 1765 14365 1777 14368
rect 1811 14396 1823 14399
rect 3050 14396 3056 14408
rect 1811 14368 3056 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3436 14405 3464 14436
rect 3881 14433 3893 14436
rect 3927 14433 3939 14467
rect 4632 14464 4660 14495
rect 5184 14464 5212 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 5629 14563 5687 14569
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8573 14603 8631 14609
rect 8573 14600 8585 14603
rect 8168 14572 8585 14600
rect 8168 14560 8174 14572
rect 8573 14569 8585 14572
rect 8619 14600 8631 14603
rect 9582 14600 9588 14612
rect 8619 14572 9588 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11517 14603 11575 14609
rect 11517 14569 11529 14603
rect 11563 14600 11575 14603
rect 11606 14600 11612 14612
rect 11563 14572 11612 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 11701 14603 11759 14609
rect 11701 14569 11713 14603
rect 11747 14600 11759 14603
rect 17310 14600 17316 14612
rect 11747 14572 17316 14600
rect 11747 14569 11759 14572
rect 11701 14563 11759 14569
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 18785 14603 18843 14609
rect 18785 14600 18797 14603
rect 18656 14572 18797 14600
rect 18656 14560 18662 14572
rect 18785 14569 18797 14572
rect 18831 14569 18843 14603
rect 18785 14563 18843 14569
rect 5258 14492 5264 14544
rect 5316 14532 5322 14544
rect 5997 14535 6055 14541
rect 5997 14532 6009 14535
rect 5316 14504 6009 14532
rect 5316 14492 5322 14504
rect 5997 14501 6009 14504
rect 6043 14501 6055 14535
rect 5997 14495 6055 14501
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14501 8815 14535
rect 11624 14532 11652 14560
rect 11974 14532 11980 14544
rect 11624 14504 11980 14532
rect 8757 14495 8815 14501
rect 3881 14427 3939 14433
rect 4356 14436 4568 14464
rect 4632 14436 4936 14464
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3602 14356 3608 14408
rect 3660 14356 3666 14408
rect 3694 14356 3700 14408
rect 3752 14396 3758 14408
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3752 14368 3801 14396
rect 3752 14356 3758 14368
rect 3789 14365 3801 14368
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 3970 14356 3976 14408
rect 4028 14356 4034 14408
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 2032 14331 2090 14337
rect 2032 14297 2044 14331
rect 2078 14328 2090 14331
rect 2130 14328 2136 14340
rect 2078 14300 2136 14328
rect 2078 14297 2090 14300
rect 2032 14291 2090 14297
rect 2130 14288 2136 14300
rect 2188 14288 2194 14340
rect 3620 14328 3648 14356
rect 4356 14328 4384 14436
rect 4433 14399 4491 14405
rect 4433 14365 4445 14399
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 3620 14300 4384 14328
rect 4448 14260 4476 14359
rect 4540 14328 4568 14436
rect 4706 14356 4712 14408
rect 4764 14356 4770 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4908 14405 4936 14436
rect 5092 14436 5212 14464
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 4982 14356 4988 14408
rect 5040 14356 5046 14408
rect 5092 14405 5120 14436
rect 5350 14424 5356 14476
rect 5408 14464 5414 14476
rect 6086 14464 6092 14476
rect 5408 14436 6092 14464
rect 5408 14424 5414 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14365 5135 14399
rect 5534 14396 5540 14408
rect 5077 14359 5135 14365
rect 5184 14368 5540 14396
rect 5092 14328 5120 14359
rect 4540 14300 5120 14328
rect 5184 14260 5212 14368
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 6236 14368 6285 14396
rect 6236 14356 6242 14368
rect 6273 14365 6285 14368
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 6546 14396 6552 14408
rect 6411 14368 6552 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 6696 14368 7113 14396
rect 6696 14356 6702 14368
rect 7101 14365 7113 14368
rect 7147 14365 7159 14399
rect 7101 14359 7159 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 8018 14396 8024 14408
rect 7423 14368 8024 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 8772 14396 8800 14495
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 17126 14492 17132 14544
rect 17184 14492 17190 14544
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 12158 14464 12164 14476
rect 11388 14436 12164 14464
rect 11388 14424 11394 14436
rect 12158 14424 12164 14436
rect 12216 14464 12222 14476
rect 12216 14436 12756 14464
rect 12216 14424 12222 14436
rect 8941 14399 8999 14405
rect 8772 14368 8892 14396
rect 5353 14331 5411 14337
rect 5353 14297 5365 14331
rect 5399 14328 5411 14331
rect 5810 14328 5816 14340
rect 5399 14300 5816 14328
rect 5399 14297 5411 14300
rect 5353 14291 5411 14297
rect 5810 14288 5816 14300
rect 5868 14288 5874 14340
rect 7561 14331 7619 14337
rect 7561 14297 7573 14331
rect 7607 14328 7619 14331
rect 8389 14331 8447 14337
rect 8389 14328 8401 14331
rect 7607 14300 8401 14328
rect 7607 14297 7619 14300
rect 7561 14291 7619 14297
rect 8389 14297 8401 14300
rect 8435 14328 8447 14331
rect 8588 14328 8616 14356
rect 8435 14300 8616 14328
rect 8864 14328 8892 14368
rect 8941 14365 8953 14399
rect 8987 14396 8999 14399
rect 9766 14396 9772 14408
rect 8987 14368 9772 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11848 14368 11897 14396
rect 11848 14356 11854 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 11974 14356 11980 14408
rect 12032 14396 12038 14408
rect 12728 14405 12756 14436
rect 12986 14424 12992 14476
rect 13044 14424 13050 14476
rect 13906 14424 13912 14476
rect 13964 14424 13970 14476
rect 18800 14464 18828 14563
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 22186 14600 22192 14612
rect 20312 14572 22192 14600
rect 20312 14560 20318 14572
rect 22186 14560 22192 14572
rect 22244 14600 22250 14612
rect 22830 14600 22836 14612
rect 22244 14572 22836 14600
rect 22244 14560 22250 14572
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 20864 14504 21680 14532
rect 20864 14492 20870 14504
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 18800 14436 19809 14464
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 21453 14467 21511 14473
rect 21453 14464 21465 14467
rect 19797 14427 19855 14433
rect 20916 14436 21465 14464
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 12032 14368 12541 14396
rect 12032 14356 12038 14368
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 15390 14399 15448 14405
rect 15390 14365 15402 14399
rect 15436 14365 15448 14399
rect 15390 14359 15448 14365
rect 9186 14331 9244 14337
rect 9186 14328 9198 14331
rect 8864 14300 9198 14328
rect 8435 14297 8447 14300
rect 8389 14291 8447 14297
rect 9186 14297 9198 14300
rect 9232 14297 9244 14331
rect 9186 14291 9244 14297
rect 11333 14331 11391 14337
rect 11333 14297 11345 14331
rect 11379 14328 11391 14331
rect 11808 14328 11836 14356
rect 11379 14300 11836 14328
rect 11379 14297 11391 14300
rect 11333 14291 11391 14297
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 15194 14328 15200 14340
rect 12676 14300 15200 14328
rect 12676 14288 12682 14300
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15405 14272 15433 14359
rect 15654 14356 15660 14408
rect 15712 14396 15718 14408
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15712 14368 15761 14396
rect 15712 14356 15718 14368
rect 15749 14365 15761 14368
rect 15795 14396 15807 14399
rect 16942 14396 16948 14408
rect 15795 14368 16948 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16942 14356 16948 14368
rect 17000 14396 17006 14408
rect 17405 14399 17463 14405
rect 17405 14396 17417 14399
rect 17000 14368 17417 14396
rect 17000 14356 17006 14368
rect 17405 14365 17417 14368
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 18506 14356 18512 14408
rect 18564 14396 18570 14408
rect 20916 14405 20944 14436
rect 21453 14433 21465 14436
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 20533 14399 20591 14405
rect 20533 14396 20545 14399
rect 18564 14368 20545 14396
rect 18564 14356 18570 14368
rect 20533 14365 20545 14368
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 20717 14359 20775 14365
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 16016 14331 16074 14337
rect 16016 14297 16028 14331
rect 16062 14328 16074 14331
rect 16666 14328 16672 14340
rect 16062 14300 16672 14328
rect 16062 14297 16074 14300
rect 16016 14291 16074 14297
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 17672 14331 17730 14337
rect 17672 14297 17684 14331
rect 17718 14328 17730 14331
rect 18598 14328 18604 14340
rect 17718 14300 18604 14328
rect 17718 14297 17730 14300
rect 17672 14291 17730 14297
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 20438 14288 20444 14340
rect 20496 14328 20502 14340
rect 20732 14328 20760 14359
rect 20496 14300 20760 14328
rect 20496 14288 20502 14300
rect 4448 14232 5212 14260
rect 5442 14220 5448 14272
rect 5500 14220 5506 14272
rect 5626 14220 5632 14272
rect 5684 14220 5690 14272
rect 6365 14263 6423 14269
rect 6365 14229 6377 14263
rect 6411 14260 6423 14263
rect 6454 14260 6460 14272
rect 6411 14232 6460 14260
rect 6411 14229 6423 14232
rect 6365 14223 6423 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7466 14260 7472 14272
rect 7239 14232 7472 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8599 14263 8657 14269
rect 8599 14229 8611 14263
rect 8645 14260 8657 14263
rect 9306 14260 9312 14272
rect 8645 14232 9312 14260
rect 8645 14229 8657 14232
rect 8599 14223 8657 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 10321 14263 10379 14269
rect 10321 14260 10333 14263
rect 9640 14232 10333 14260
rect 9640 14220 9646 14232
rect 10321 14229 10333 14232
rect 10367 14229 10379 14263
rect 10321 14223 10379 14229
rect 11543 14263 11601 14269
rect 11543 14229 11555 14263
rect 11589 14260 11601 14263
rect 12342 14260 12348 14272
rect 11589 14232 12348 14260
rect 11589 14229 11601 14232
rect 11543 14223 11601 14229
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14260 13323 14263
rect 13538 14260 13544 14272
rect 13311 14232 13544 14260
rect 13311 14229 13323 14232
rect 13265 14223 13323 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 15286 14260 15292 14272
rect 14323 14232 15292 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 15378 14220 15384 14272
rect 15436 14220 15442 14272
rect 18966 14220 18972 14272
rect 19024 14260 19030 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 19024 14232 19257 14260
rect 19024 14220 19030 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19852 14232 19993 14260
rect 19852 14220 19858 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21008 14260 21036 14359
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 21652 14405 21680 14504
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 23382 14396 23388 14408
rect 21683 14368 23388 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 23382 14356 23388 14368
rect 23440 14356 23446 14408
rect 24394 14356 24400 14408
rect 24452 14356 24458 14408
rect 21100 14328 21128 14356
rect 21100 14300 21772 14328
rect 20772 14232 21036 14260
rect 20772 14220 20778 14232
rect 21358 14220 21364 14272
rect 21416 14220 21422 14272
rect 21744 14260 21772 14300
rect 21818 14288 21824 14340
rect 21876 14288 21882 14340
rect 24302 14288 24308 14340
rect 24360 14328 24366 14340
rect 24642 14331 24700 14337
rect 24642 14328 24654 14331
rect 24360 14300 24654 14328
rect 24360 14288 24366 14300
rect 24642 14297 24654 14300
rect 24688 14297 24700 14331
rect 24642 14291 24700 14297
rect 23198 14260 23204 14272
rect 21744 14232 23204 14260
rect 23198 14220 23204 14232
rect 23256 14260 23262 14272
rect 24026 14260 24032 14272
rect 23256 14232 24032 14260
rect 23256 14220 23262 14232
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 25777 14263 25835 14269
rect 25777 14260 25789 14263
rect 25740 14232 25789 14260
rect 25740 14220 25746 14232
rect 25777 14229 25789 14232
rect 25823 14229 25835 14263
rect 25777 14223 25835 14229
rect 1104 14170 26220 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 26220 14170
rect 1104 14096 26220 14118
rect 106 14016 112 14068
rect 164 14056 170 14068
rect 164 14028 13308 14056
rect 164 14016 170 14028
rect 3145 13991 3203 13997
rect 3145 13957 3157 13991
rect 3191 13988 3203 13991
rect 3191 13960 3372 13988
rect 3191 13957 3203 13960
rect 3145 13951 3203 13957
rect 1578 13880 1584 13932
rect 1636 13880 1642 13932
rect 1854 13929 1860 13932
rect 1848 13920 1860 13929
rect 1815 13892 1860 13920
rect 1848 13883 1860 13892
rect 1854 13880 1860 13883
rect 1912 13880 1918 13932
rect 2958 13880 2964 13932
rect 3016 13920 3022 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 3016 13892 3065 13920
rect 3016 13880 3022 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 3234 13880 3240 13932
rect 3292 13880 3298 13932
rect 3344 13929 3372 13960
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 5721 13991 5779 13997
rect 5316 13960 5488 13988
rect 5316 13948 5322 13960
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 3786 13920 3792 13932
rect 3559 13892 3792 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 2924 13824 3004 13852
rect 2924 13812 2930 13824
rect 2976 13793 3004 13824
rect 3142 13812 3148 13864
rect 3200 13852 3206 13864
rect 3528 13852 3556 13883
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4856 13892 4905 13920
rect 4856 13880 4862 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13889 5227 13923
rect 5169 13883 5227 13889
rect 3200 13824 3556 13852
rect 3200 13812 3206 13824
rect 2961 13787 3019 13793
rect 2961 13753 2973 13787
rect 3007 13753 3019 13787
rect 2961 13747 3019 13753
rect 3326 13676 3332 13728
rect 3384 13676 3390 13728
rect 4982 13676 4988 13728
rect 5040 13676 5046 13728
rect 5184 13716 5212 13883
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5460 13929 5488 13960
rect 5721 13957 5733 13991
rect 5767 13988 5779 13991
rect 6270 13988 6276 14000
rect 5767 13960 6276 13988
rect 5767 13957 5779 13960
rect 5721 13951 5779 13957
rect 6270 13948 6276 13960
rect 6328 13988 6334 14000
rect 6365 13991 6423 13997
rect 6365 13988 6377 13991
rect 6328 13960 6377 13988
rect 6328 13948 6334 13960
rect 6365 13957 6377 13960
rect 6411 13957 6423 13991
rect 6365 13951 6423 13957
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6565 13991 6623 13997
rect 6565 13988 6577 13991
rect 6512 13960 6577 13988
rect 6512 13948 6518 13960
rect 6565 13957 6577 13960
rect 6611 13957 6623 13991
rect 6565 13951 6623 13957
rect 6656 13960 7788 13988
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 5810 13880 5816 13932
rect 5868 13880 5874 13932
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13889 5963 13923
rect 5905 13883 5963 13889
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5920 13852 5948 13883
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6656 13920 6684 13960
rect 7760 13932 7788 13960
rect 8018 13948 8024 14000
rect 8076 13948 8082 14000
rect 8294 13948 8300 14000
rect 8352 13948 8358 14000
rect 8754 13988 8760 14000
rect 8588 13960 8760 13988
rect 8296 13945 8354 13948
rect 7101 13923 7159 13929
rect 7101 13920 7113 13923
rect 6052 13892 6684 13920
rect 6748 13892 7113 13920
rect 6052 13880 6058 13892
rect 6638 13852 6644 13864
rect 5307 13824 5948 13852
rect 6104 13824 6644 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 5626 13784 5632 13796
rect 5408 13756 5632 13784
rect 5408 13744 5414 13756
rect 5626 13744 5632 13756
rect 5684 13744 5690 13796
rect 5994 13784 6000 13796
rect 5736 13756 6000 13784
rect 5736 13716 5764 13756
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 6104 13793 6132 13824
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 6748 13793 6776 13892
rect 7101 13889 7113 13892
rect 7147 13889 7159 13923
rect 7101 13883 7159 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7466 13920 7472 13932
rect 7423 13892 7472 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7800 13892 8248 13920
rect 8296 13911 8308 13945
rect 8342 13911 8354 13945
rect 8588 13929 8616 13960
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 9398 13948 9404 14000
rect 9456 13948 9462 14000
rect 9490 13948 9496 14000
rect 9548 13988 9554 14000
rect 9601 13991 9659 13997
rect 9601 13988 9613 13991
rect 9548 13960 9613 13988
rect 9548 13948 9554 13960
rect 9601 13957 9613 13960
rect 9647 13957 9659 13991
rect 9953 13991 10011 13997
rect 9953 13988 9965 13991
rect 9601 13951 9659 13957
rect 9692 13960 9965 13988
rect 8296 13905 8354 13911
rect 8389 13921 8447 13927
rect 7800 13880 7806 13892
rect 8018 13812 8024 13864
rect 8076 13812 8082 13864
rect 6089 13787 6147 13793
rect 6089 13753 6101 13787
rect 6135 13753 6147 13787
rect 6089 13747 6147 13753
rect 6733 13787 6791 13793
rect 6733 13753 6745 13787
rect 6779 13753 6791 13787
rect 6733 13747 6791 13753
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 8110 13784 8116 13796
rect 7340 13756 8116 13784
rect 7340 13744 7346 13756
rect 8110 13744 8116 13756
rect 8168 13744 8174 13796
rect 8220 13784 8248 13892
rect 8389 13887 8401 13921
rect 8435 13887 8447 13921
rect 8389 13881 8447 13887
rect 8573 13923 8631 13929
rect 8573 13889 8585 13923
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 8671 13923 8729 13929
rect 8671 13889 8683 13923
rect 8717 13889 8729 13923
rect 8671 13883 8729 13889
rect 8404 13852 8432 13881
rect 8478 13852 8484 13864
rect 8404 13824 8484 13852
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8588 13784 8616 13883
rect 8686 13852 8714 13883
rect 8846 13880 8852 13932
rect 8904 13880 8910 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9033 13923 9091 13929
rect 8987 13889 9000 13920
rect 8941 13883 9000 13889
rect 9033 13889 9045 13923
rect 9079 13918 9091 13923
rect 9122 13918 9128 13932
rect 9079 13890 9128 13918
rect 9079 13889 9091 13890
rect 9033 13883 9091 13889
rect 8686 13824 8717 13852
rect 8220 13756 8616 13784
rect 5184 13688 5764 13716
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 5868 13688 6561 13716
rect 5868 13676 5874 13688
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 6549 13679 6607 13685
rect 7834 13676 7840 13728
rect 7892 13716 7898 13728
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7892 13688 8217 13716
rect 7892 13676 7898 13688
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 8205 13679 8263 13685
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8352 13688 8493 13716
rect 8352 13676 8358 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8689 13716 8717 13824
rect 8972 13844 9000 13883
rect 9122 13880 9128 13890
rect 9180 13880 9186 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9692 13920 9720 13960
rect 9953 13957 9965 13960
rect 9999 13957 10011 13991
rect 9953 13951 10011 13957
rect 12158 13948 12164 14000
rect 12216 13948 12222 14000
rect 13280 13997 13308 14028
rect 14734 14016 14740 14068
rect 14792 14016 14798 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 16206 14056 16212 14068
rect 15896 14028 16212 14056
rect 15896 14016 15902 14028
rect 16206 14016 16212 14028
rect 16264 14056 16270 14068
rect 16485 14059 16543 14065
rect 16485 14056 16497 14059
rect 16264 14028 16497 14056
rect 16264 14016 16270 14028
rect 16485 14025 16497 14028
rect 16531 14025 16543 14059
rect 16485 14019 16543 14025
rect 18506 14016 18512 14068
rect 18564 14016 18570 14068
rect 18598 14016 18604 14068
rect 18656 14016 18662 14068
rect 18966 14016 18972 14068
rect 19024 14016 19030 14068
rect 19429 14059 19487 14065
rect 19429 14025 19441 14059
rect 19475 14025 19487 14059
rect 19429 14019 19487 14025
rect 15378 13997 15384 14000
rect 12437 13991 12495 13997
rect 12437 13957 12449 13991
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 12653 13991 12711 13997
rect 12653 13957 12665 13991
rect 12699 13988 12711 13991
rect 12989 13991 13047 13997
rect 12989 13988 13001 13991
rect 12699 13960 13001 13988
rect 12699 13957 12711 13960
rect 12653 13951 12711 13957
rect 12989 13957 13001 13960
rect 13035 13957 13047 13991
rect 12989 13951 13047 13957
rect 13265 13991 13323 13997
rect 13265 13957 13277 13991
rect 13311 13957 13323 13991
rect 13265 13951 13323 13957
rect 15350 13991 15384 13997
rect 15350 13957 15362 13991
rect 15350 13951 15384 13957
rect 9364 13892 9720 13920
rect 9861 13923 9919 13929
rect 9364 13880 9370 13892
rect 9861 13889 9873 13923
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 9876 13852 9904 13883
rect 10042 13880 10048 13932
rect 10100 13880 10106 13932
rect 11790 13880 11796 13932
rect 11848 13880 11854 13932
rect 12452 13920 12480 13951
rect 15378 13948 15384 13951
rect 15436 13948 15442 14000
rect 17396 13991 17454 13997
rect 17396 13957 17408 13991
rect 17442 13988 17454 13991
rect 19444 13988 19472 14019
rect 19794 14016 19800 14068
rect 19852 14016 19858 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 21082 14056 21088 14068
rect 20128 14028 21088 14056
rect 20128 14016 20134 14028
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21358 14016 21364 14068
rect 21416 14056 21422 14068
rect 23201 14059 23259 14065
rect 21416 14028 22094 14056
rect 21416 14016 21422 14028
rect 22066 13997 22094 14028
rect 23201 14025 23213 14059
rect 23247 14056 23259 14059
rect 23382 14056 23388 14068
rect 23247 14028 23388 14056
rect 23247 14025 23259 14028
rect 23201 14019 23259 14025
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 24302 14016 24308 14068
rect 24360 14016 24366 14068
rect 25406 14016 25412 14068
rect 25464 14016 25470 14068
rect 25774 14016 25780 14068
rect 25832 14016 25838 14068
rect 22066 13991 22124 13997
rect 17442 13960 19472 13988
rect 20272 13960 20944 13988
rect 17442 13957 17454 13960
rect 17396 13951 17454 13957
rect 12802 13920 12808 13932
rect 12452 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13078 13880 13084 13932
rect 13136 13880 13142 13932
rect 15102 13880 15108 13932
rect 15160 13880 15166 13932
rect 16850 13920 16856 13932
rect 15212 13892 16856 13920
rect 12618 13852 12624 13864
rect 9201 13844 9904 13852
rect 8972 13824 9904 13844
rect 12360 13824 12624 13852
rect 8972 13816 9229 13824
rect 9784 13793 9812 13824
rect 12360 13793 12388 13824
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 13630 13852 13636 13864
rect 12820 13824 13636 13852
rect 12820 13793 12848 13824
rect 13630 13812 13636 13824
rect 13688 13852 13694 13864
rect 15212 13852 15240 13892
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17129 13923 17187 13929
rect 17129 13920 17141 13923
rect 17000 13892 17141 13920
rect 17000 13880 17006 13892
rect 17129 13889 17141 13892
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13920 19119 13923
rect 19518 13920 19524 13932
rect 19107 13892 19524 13920
rect 19107 13889 19119 13892
rect 19061 13883 19119 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20162 13920 20168 13932
rect 19935 13892 20168 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20272 13929 20300 13960
rect 20916 13932 20944 13960
rect 22066 13957 22078 13991
rect 22112 13957 22124 13991
rect 22066 13951 22124 13957
rect 23750 13948 23756 14000
rect 23808 13988 23814 14000
rect 24486 13988 24492 14000
rect 23808 13960 23980 13988
rect 23808 13948 23814 13960
rect 20257 13923 20315 13929
rect 20257 13889 20269 13923
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20513 13923 20571 13929
rect 20513 13920 20525 13923
rect 20404 13892 20525 13920
rect 20404 13880 20410 13892
rect 20513 13889 20525 13892
rect 20559 13889 20571 13923
rect 20513 13883 20571 13889
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 21634 13920 21640 13932
rect 20956 13892 21640 13920
rect 20956 13880 20962 13892
rect 21634 13880 21640 13892
rect 21692 13920 21698 13932
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21692 13892 21833 13920
rect 21692 13880 21698 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 21910 13880 21916 13932
rect 21968 13880 21974 13932
rect 23952 13929 23980 13960
rect 24044 13960 24492 13988
rect 24044 13932 24072 13960
rect 24486 13948 24492 13960
rect 24544 13948 24550 14000
rect 24581 13991 24639 13997
rect 24581 13957 24593 13991
rect 24627 13988 24639 13991
rect 25682 13988 25688 14000
rect 24627 13960 25688 13988
rect 24627 13957 24639 13960
rect 24581 13951 24639 13957
rect 25682 13948 25688 13960
rect 25740 13948 25746 14000
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13889 23903 13923
rect 23845 13883 23903 13889
rect 23937 13923 23995 13929
rect 23937 13889 23949 13923
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 13688 13824 15240 13852
rect 19153 13855 19211 13861
rect 13688 13812 13694 13824
rect 19153 13821 19165 13855
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13821 20039 13855
rect 21928 13852 21956 13880
rect 19981 13815 20039 13821
rect 21376 13824 21956 13852
rect 9769 13787 9827 13793
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 12345 13787 12403 13793
rect 9815 13756 9849 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 12345 13753 12357 13787
rect 12391 13753 12403 13787
rect 12345 13747 12403 13753
rect 12805 13787 12863 13793
rect 12805 13753 12817 13787
rect 12851 13753 12863 13787
rect 12805 13747 12863 13753
rect 18322 13744 18328 13796
rect 18380 13784 18386 13796
rect 19168 13784 19196 13815
rect 19996 13784 20024 13815
rect 18380 13756 20024 13784
rect 18380 13744 18386 13756
rect 9030 13716 9036 13728
rect 8689 13688 9036 13716
rect 8481 13679 8539 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 9272 13688 9321 13716
rect 9272 13676 9278 13688
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 9582 13676 9588 13728
rect 9640 13676 9646 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12066 13716 12072 13728
rect 11940 13688 12072 13716
rect 11940 13676 11946 13688
rect 12066 13676 12072 13688
rect 12124 13716 12130 13728
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 12124 13688 12173 13716
rect 12124 13676 12130 13688
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 12161 13679 12219 13685
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12492 13688 12633 13716
rect 12492 13676 12498 13688
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 12621 13679 12679 13685
rect 20438 13676 20444 13728
rect 20496 13716 20502 13728
rect 21376 13716 21404 13824
rect 21450 13744 21456 13796
rect 21508 13784 21514 13796
rect 21637 13787 21695 13793
rect 21637 13784 21649 13787
rect 21508 13756 21649 13784
rect 21508 13744 21514 13756
rect 21637 13753 21649 13756
rect 21683 13784 21695 13787
rect 21726 13784 21732 13796
rect 21683 13756 21732 13784
rect 21683 13753 21695 13756
rect 21637 13747 21695 13753
rect 21726 13744 21732 13756
rect 21784 13744 21790 13796
rect 23676 13784 23704 13883
rect 23860 13852 23888 13883
rect 24026 13880 24032 13932
rect 24084 13880 24090 13932
rect 24118 13880 24124 13932
rect 24176 13920 24182 13932
rect 24397 13923 24455 13929
rect 24397 13920 24409 13923
rect 24176 13892 24409 13920
rect 24176 13880 24182 13892
rect 24397 13889 24409 13892
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 24765 13855 24823 13861
rect 24765 13852 24777 13855
rect 23860 13824 24777 13852
rect 24765 13821 24777 13824
rect 24811 13821 24823 13855
rect 24765 13815 24823 13821
rect 22848 13756 23704 13784
rect 20496 13688 21404 13716
rect 20496 13676 20502 13688
rect 21542 13676 21548 13728
rect 21600 13716 21606 13728
rect 22848 13716 22876 13756
rect 21600 13688 22876 13716
rect 21600 13676 21606 13688
rect 22922 13676 22928 13728
rect 22980 13716 22986 13728
rect 25608 13716 25636 13883
rect 22980 13688 25636 13716
rect 22980 13676 22986 13688
rect 1104 13626 26220 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 26220 13626
rect 1104 13552 26220 13574
rect 2130 13472 2136 13524
rect 2188 13472 2194 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2590 13512 2596 13524
rect 2363 13484 2596 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5258 13512 5264 13524
rect 5215 13484 5264 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 6270 13472 6276 13524
rect 6328 13472 6334 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 7064 13484 7113 13512
rect 7064 13472 7070 13484
rect 7101 13481 7113 13484
rect 7147 13481 7159 13515
rect 7101 13475 7159 13481
rect 7466 13472 7472 13524
rect 7524 13472 7530 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 8076 13484 8217 13512
rect 8076 13472 8082 13484
rect 8205 13481 8217 13484
rect 8251 13481 8263 13515
rect 8205 13475 8263 13481
rect 8665 13515 8723 13521
rect 8665 13481 8677 13515
rect 8711 13512 8723 13515
rect 8754 13512 8760 13524
rect 8711 13484 8760 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 10042 13512 10048 13524
rect 9263 13484 10048 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 13998 13512 14004 13524
rect 13955 13484 14004 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15436 13484 15577 13512
rect 15436 13472 15442 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 18230 13472 18236 13524
rect 18288 13512 18294 13524
rect 18509 13515 18567 13521
rect 18509 13512 18521 13515
rect 18288 13484 18521 13512
rect 18288 13472 18294 13484
rect 18509 13481 18521 13484
rect 18555 13481 18567 13515
rect 18509 13475 18567 13481
rect 20165 13515 20223 13521
rect 20165 13481 20177 13515
rect 20211 13512 20223 13515
rect 20346 13512 20352 13524
rect 20211 13484 20352 13512
rect 20211 13481 20223 13484
rect 20165 13475 20223 13481
rect 5442 13404 5448 13456
rect 5500 13404 5506 13456
rect 5537 13447 5595 13453
rect 5537 13413 5549 13447
rect 5583 13444 5595 13447
rect 6178 13444 6184 13456
rect 5583 13416 6184 13444
rect 5583 13413 5595 13416
rect 5537 13407 5595 13413
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 6917 13447 6975 13453
rect 6917 13413 6929 13447
rect 6963 13444 6975 13447
rect 6963 13416 8432 13444
rect 6963 13413 6975 13416
rect 6917 13407 6975 13413
rect 7628 13379 7686 13385
rect 5644 13348 6132 13376
rect 5644 13320 5672 13348
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5040 13280 5365 13308
rect 5040 13268 5046 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 6104 13317 6132 13348
rect 7628 13345 7640 13379
rect 7674 13376 7686 13379
rect 8294 13376 8300 13388
rect 7674 13348 8300 13376
rect 7674 13345 7686 13348
rect 7628 13339 7686 13345
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5776 13280 5825 13308
rect 5776 13268 5782 13280
rect 5813 13277 5825 13280
rect 5859 13308 5871 13311
rect 5905 13311 5963 13317
rect 5905 13308 5917 13311
rect 5859 13280 5917 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 5905 13277 5917 13280
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6880 13280 7113 13308
rect 6880 13268 6886 13280
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 2501 13243 2559 13249
rect 2501 13209 2513 13243
rect 2547 13240 2559 13243
rect 2682 13240 2688 13252
rect 2547 13212 2688 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 2682 13200 2688 13212
rect 2740 13200 2746 13252
rect 2301 13175 2359 13181
rect 2301 13141 2313 13175
rect 2347 13172 2359 13175
rect 3326 13172 3332 13184
rect 2347 13144 3332 13172
rect 2347 13141 2359 13144
rect 2301 13135 2359 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 7208 13172 7236 13271
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7745 13311 7803 13317
rect 7745 13308 7757 13311
rect 7524 13280 7757 13308
rect 7524 13268 7530 13280
rect 7745 13277 7757 13280
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 7834 13268 7840 13320
rect 7892 13268 7898 13320
rect 8110 13308 8116 13320
rect 7944 13280 8116 13308
rect 7377 13243 7435 13249
rect 7377 13209 7389 13243
rect 7423 13240 7435 13243
rect 7944 13240 7972 13280
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8404 13317 8432 13416
rect 9122 13376 9128 13388
rect 8772 13348 9128 13376
rect 8772 13317 8800 13348
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 14921 13379 14979 13385
rect 14921 13376 14933 13379
rect 13412 13348 14933 13376
rect 13412 13336 13418 13348
rect 14921 13345 14933 13348
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8481 13271 8539 13277
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13308 8999 13311
rect 9490 13308 9496 13320
rect 8987 13280 9496 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 7423 13212 7972 13240
rect 7423 13209 7435 13212
rect 7377 13203 7435 13209
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8496 13240 8524 13271
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 8260 13212 8524 13240
rect 8260 13200 8266 13212
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9217 13243 9275 13249
rect 9217 13240 9229 13243
rect 8720 13212 9229 13240
rect 8720 13200 8726 13212
rect 9217 13209 9229 13212
rect 9263 13240 9275 13243
rect 9582 13240 9588 13252
rect 9263 13212 9588 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 12268 13240 12296 13271
rect 12434 13268 12440 13320
rect 12492 13268 12498 13320
rect 13538 13268 13544 13320
rect 13596 13268 13602 13320
rect 14936 13308 14964 13339
rect 16206 13336 16212 13388
rect 16264 13336 16270 13388
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 17000 13348 17141 13376
rect 17000 13336 17006 13348
rect 17129 13345 17141 13348
rect 17175 13345 17187 13379
rect 18524 13376 18552 13475
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 20806 13472 20812 13524
rect 20864 13472 20870 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21542 13512 21548 13524
rect 21140 13484 21548 13512
rect 21140 13472 21146 13484
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 21910 13472 21916 13524
rect 21968 13512 21974 13524
rect 21968 13484 22094 13512
rect 21968 13472 21974 13484
rect 19886 13404 19892 13456
rect 19944 13444 19950 13456
rect 20824 13444 20852 13472
rect 19944 13416 20852 13444
rect 19944 13404 19950 13416
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 18524 13348 19809 13376
rect 17129 13339 17187 13345
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 20898 13336 20904 13388
rect 20956 13336 20962 13388
rect 18230 13308 18236 13320
rect 14936 13280 18236 13308
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 20254 13268 20260 13320
rect 20312 13308 20318 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 20312 13280 20453 13308
rect 20312 13268 20318 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21542 13308 21548 13320
rect 20855 13280 21548 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 12986 13240 12992 13252
rect 12268 13212 12992 13240
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 13449 13243 13507 13249
rect 13449 13209 13461 13243
rect 13495 13240 13507 13243
rect 14274 13240 14280 13252
rect 13495 13212 14280 13240
rect 13495 13209 13507 13212
rect 13449 13203 13507 13209
rect 14274 13200 14280 13212
rect 14332 13200 14338 13252
rect 15105 13243 15163 13249
rect 15105 13209 15117 13243
rect 15151 13240 15163 13243
rect 15286 13240 15292 13252
rect 15151 13212 15292 13240
rect 15151 13209 15163 13212
rect 15105 13203 15163 13209
rect 15286 13200 15292 13212
rect 15344 13200 15350 13252
rect 17396 13243 17454 13249
rect 17396 13209 17408 13243
rect 17442 13240 17454 13243
rect 17862 13240 17868 13252
rect 17442 13212 17868 13240
rect 17442 13209 17454 13212
rect 17396 13203 17454 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 8018 13172 8024 13184
rect 7208 13144 8024 13172
rect 8018 13132 8024 13144
rect 8076 13172 8082 13184
rect 8478 13172 8484 13184
rect 8076 13144 8484 13172
rect 8076 13132 8082 13144
rect 8478 13132 8484 13144
rect 8536 13172 8542 13184
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8536 13144 9045 13172
rect 8536 13132 8542 13144
rect 9033 13141 9045 13144
rect 9079 13172 9091 13175
rect 9306 13172 9312 13184
rect 9079 13144 9312 13172
rect 9079 13141 9091 13144
rect 9033 13135 9091 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 12066 13132 12072 13184
rect 12124 13132 12130 13184
rect 15197 13175 15255 13181
rect 15197 13141 15209 13175
rect 15243 13172 15255 13175
rect 15657 13175 15715 13181
rect 15657 13172 15669 13175
rect 15243 13144 15669 13172
rect 15243 13141 15255 13144
rect 15197 13135 15255 13141
rect 15657 13141 15669 13144
rect 15703 13141 15715 13175
rect 15657 13135 15715 13141
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 20640 13172 20668 13271
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22066 13308 22094 13484
rect 23198 13404 23204 13456
rect 23256 13444 23262 13456
rect 24118 13444 24124 13456
rect 23256 13416 24124 13444
rect 23256 13404 23262 13416
rect 24118 13404 24124 13416
rect 24176 13404 24182 13456
rect 23477 13379 23535 13385
rect 23477 13345 23489 13379
rect 23523 13376 23535 13379
rect 23523 13348 23796 13376
rect 23523 13345 23535 13348
rect 23477 13339 23535 13345
rect 23382 13308 23388 13320
rect 22066 13280 23388 13308
rect 23382 13268 23388 13280
rect 23440 13308 23446 13320
rect 23768 13317 23796 13348
rect 23569 13311 23627 13317
rect 23569 13308 23581 13311
rect 23440 13280 23581 13308
rect 23440 13268 23446 13280
rect 23569 13277 23581 13280
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 23753 13311 23811 13317
rect 23753 13277 23765 13311
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 21174 13249 21180 13252
rect 21168 13203 21180 13249
rect 21174 13200 21180 13203
rect 21232 13200 21238 13252
rect 21818 13200 21824 13252
rect 21876 13240 21882 13252
rect 22373 13243 22431 13249
rect 22373 13240 22385 13243
rect 21876 13212 22385 13240
rect 21876 13200 21882 13212
rect 22373 13209 22385 13212
rect 22419 13209 22431 13243
rect 22373 13203 22431 13209
rect 22557 13243 22615 13249
rect 22557 13209 22569 13243
rect 22603 13240 22615 13243
rect 22922 13240 22928 13252
rect 22603 13212 22928 13240
rect 22603 13209 22615 13212
rect 22557 13203 22615 13209
rect 21266 13172 21272 13184
rect 20640 13144 21272 13172
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22281 13175 22339 13181
rect 22281 13172 22293 13175
rect 22152 13144 22293 13172
rect 22152 13132 22158 13144
rect 22281 13141 22293 13144
rect 22327 13172 22339 13175
rect 22572 13172 22600 13203
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 23109 13243 23167 13249
rect 23109 13209 23121 13243
rect 23155 13240 23167 13243
rect 23198 13240 23204 13252
rect 23155 13212 23204 13240
rect 23155 13209 23167 13212
rect 23109 13203 23167 13209
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 23293 13243 23351 13249
rect 23293 13209 23305 13243
rect 23339 13209 23351 13243
rect 23293 13203 23351 13209
rect 22327 13144 22600 13172
rect 22327 13141 22339 13144
rect 22281 13135 22339 13141
rect 22738 13132 22744 13184
rect 22796 13132 22802 13184
rect 23308 13172 23336 13203
rect 23658 13200 23664 13252
rect 23716 13240 23722 13252
rect 23860 13240 23888 13271
rect 23934 13268 23940 13320
rect 23992 13268 23998 13320
rect 24026 13268 24032 13320
rect 24084 13308 24090 13320
rect 24394 13308 24400 13320
rect 24084 13280 24400 13308
rect 24084 13268 24090 13280
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 23716 13212 23888 13240
rect 23952 13240 23980 13268
rect 24118 13240 24124 13252
rect 23952 13212 24124 13240
rect 23716 13200 23722 13212
rect 24118 13200 24124 13212
rect 24176 13200 24182 13252
rect 24213 13243 24271 13249
rect 24213 13209 24225 13243
rect 24259 13240 24271 13243
rect 24642 13243 24700 13249
rect 24642 13240 24654 13243
rect 24259 13212 24654 13240
rect 24259 13209 24271 13212
rect 24213 13203 24271 13209
rect 24642 13209 24654 13212
rect 24688 13209 24700 13243
rect 24642 13203 24700 13209
rect 23934 13172 23940 13184
rect 23308 13144 23940 13172
rect 23934 13132 23940 13144
rect 23992 13172 23998 13184
rect 25590 13172 25596 13184
rect 23992 13144 25596 13172
rect 23992 13132 23998 13144
rect 25590 13132 25596 13144
rect 25648 13172 25654 13184
rect 25777 13175 25835 13181
rect 25777 13172 25789 13175
rect 25648 13144 25789 13172
rect 25648 13132 25654 13144
rect 25777 13141 25789 13144
rect 25823 13141 25835 13175
rect 25777 13135 25835 13141
rect 1104 13082 26220 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 26220 13082
rect 1104 13008 26220 13030
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 6178 12968 6184 12980
rect 5123 12940 6184 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 8021 12971 8079 12977
rect 8021 12968 8033 12971
rect 7892 12940 8033 12968
rect 7892 12928 7898 12940
rect 8021 12937 8033 12940
rect 8067 12937 8079 12971
rect 8021 12931 8079 12937
rect 8110 12928 8116 12980
rect 8168 12928 8174 12980
rect 8386 12968 8392 12980
rect 8312 12940 8392 12968
rect 5537 12903 5595 12909
rect 5537 12869 5549 12903
rect 5583 12900 5595 12903
rect 5810 12900 5816 12912
rect 5583 12872 5816 12900
rect 5583 12869 5595 12872
rect 5537 12863 5595 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 7653 12903 7711 12909
rect 7653 12869 7665 12903
rect 7699 12900 7711 12903
rect 7742 12900 7748 12912
rect 7699 12872 7748 12900
rect 7699 12869 7711 12872
rect 7653 12863 7711 12869
rect 7742 12860 7748 12872
rect 7800 12860 7806 12912
rect 8312 12909 8340 12940
rect 8386 12928 8392 12940
rect 8444 12968 8450 12980
rect 8662 12968 8668 12980
rect 8444 12940 8668 12968
rect 8444 12928 8450 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9125 12971 9183 12977
rect 9125 12937 9137 12971
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 8297 12903 8355 12909
rect 8297 12869 8309 12903
rect 8343 12869 8355 12903
rect 8297 12863 8355 12869
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 8628 12872 8769 12900
rect 8628 12860 8634 12872
rect 8757 12869 8769 12872
rect 8803 12869 8815 12903
rect 8757 12863 8815 12869
rect 8938 12860 8944 12912
rect 8996 12909 9002 12912
rect 8996 12903 9015 12909
rect 9003 12869 9015 12903
rect 9140 12900 9168 12931
rect 17862 12928 17868 12980
rect 17920 12928 17926 12980
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 19242 12968 19248 12980
rect 18279 12940 19248 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19518 12928 19524 12980
rect 19576 12928 19582 12980
rect 21174 12928 21180 12980
rect 21232 12928 21238 12980
rect 21266 12928 21272 12980
rect 21324 12928 21330 12980
rect 24118 12968 24124 12980
rect 23400 12940 24124 12968
rect 10330 12903 10388 12909
rect 10330 12900 10342 12903
rect 9140 12872 10342 12900
rect 8996 12863 9015 12869
rect 10330 12869 10342 12872
rect 10376 12869 10388 12903
rect 22738 12900 22744 12912
rect 10330 12863 10388 12869
rect 19996 12872 20668 12900
rect 8996 12860 9002 12863
rect 2866 12792 2872 12844
rect 2924 12792 2930 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 4614 12832 4620 12844
rect 3099 12804 4620 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 4856 12736 5089 12764
rect 4856 12724 4862 12736
rect 5077 12733 5089 12736
rect 5123 12733 5135 12767
rect 5368 12764 5396 12795
rect 5442 12792 5448 12844
rect 5500 12792 5506 12844
rect 5718 12792 5724 12844
rect 5776 12792 5782 12844
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8018 12832 8024 12844
rect 7883 12804 8024 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 11968 12835 12026 12841
rect 11968 12801 11980 12835
rect 12014 12832 12026 12835
rect 12894 12832 12900 12844
rect 12014 12804 12900 12832
rect 12014 12801 12026 12804
rect 11968 12795 12026 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12832 18383 12835
rect 19610 12832 19616 12844
rect 18371 12804 19616 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 19886 12832 19892 12844
rect 19843 12804 19892 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 19996 12841 20024 12872
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 6822 12764 6828 12776
rect 5368 12736 6828 12764
rect 5077 12727 5135 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 10597 12767 10655 12773
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10962 12764 10968 12776
rect 10643 12736 10968 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10962 12724 10968 12736
rect 11020 12764 11026 12776
rect 11701 12767 11759 12773
rect 11701 12764 11713 12767
rect 11020 12736 11713 12764
rect 11020 12724 11026 12736
rect 11701 12733 11713 12736
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 18288 12736 18429 12764
rect 18288 12724 18294 12736
rect 18417 12733 18429 12736
rect 18463 12764 18475 12767
rect 19058 12764 19064 12776
rect 18463 12736 19064 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 20088 12764 20116 12795
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 20496 12804 20545 12832
rect 20496 12792 20502 12804
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 19576 12736 20116 12764
rect 19576 12724 19582 12736
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 5592 12668 5733 12696
rect 5592 12656 5598 12668
rect 5721 12665 5733 12668
rect 5767 12665 5779 12699
rect 20640 12696 20668 12872
rect 20732 12872 22744 12900
rect 20732 12841 20760 12872
rect 22738 12860 22744 12872
rect 22796 12860 22802 12912
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 20806 12792 20812 12844
rect 20864 12792 20870 12844
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12832 20959 12835
rect 21174 12832 21180 12844
rect 20947 12804 21180 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 21634 12792 21640 12844
rect 21692 12792 21698 12844
rect 23400 12832 23428 12940
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 25774 12928 25780 12980
rect 25832 12928 25838 12980
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 23753 12903 23811 12909
rect 23753 12900 23765 12903
rect 23532 12872 23765 12900
rect 23532 12860 23538 12872
rect 23753 12869 23765 12872
rect 23799 12869 23811 12903
rect 23753 12863 23811 12869
rect 21744 12804 23428 12832
rect 21192 12764 21220 12792
rect 21744 12764 21772 12804
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 23658 12792 23664 12844
rect 23716 12792 23722 12844
rect 23934 12792 23940 12844
rect 23992 12792 23998 12844
rect 24026 12792 24032 12844
rect 24084 12792 24090 12844
rect 24296 12835 24354 12841
rect 24296 12801 24308 12835
rect 24342 12832 24354 12835
rect 25038 12832 25044 12844
rect 24342 12804 25044 12832
rect 24342 12801 24354 12804
rect 24296 12795 24354 12801
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25590 12792 25596 12844
rect 25648 12841 25654 12844
rect 25648 12832 25657 12841
rect 25648 12804 25693 12832
rect 25648 12795 25657 12804
rect 25648 12792 25654 12795
rect 21192 12736 21772 12764
rect 22002 12724 22008 12776
rect 22060 12764 22066 12776
rect 23750 12764 23756 12776
rect 22060 12736 23756 12764
rect 22060 12724 22066 12736
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 20640 12668 23612 12696
rect 5721 12659 5779 12665
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3418 12628 3424 12640
rect 3099 12600 3424 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4764 12600 5273 12628
rect 4764 12588 4770 12600
rect 5261 12597 5273 12600
rect 5307 12597 5319 12631
rect 5261 12591 5319 12597
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 8941 12631 8999 12637
rect 8941 12628 8953 12631
rect 7340 12600 8953 12628
rect 7340 12588 7346 12600
rect 8941 12597 8953 12600
rect 8987 12597 8999 12631
rect 8941 12591 8999 12597
rect 9217 12631 9275 12637
rect 9217 12597 9229 12631
rect 9263 12628 9275 12631
rect 9306 12628 9312 12640
rect 9263 12600 9312 12628
rect 9263 12597 9275 12600
rect 9217 12591 9275 12597
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 13081 12631 13139 12637
rect 13081 12597 13093 12631
rect 13127 12628 13139 12631
rect 13262 12628 13268 12640
rect 13127 12600 13268 12628
rect 13127 12597 13139 12600
rect 13081 12591 13139 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 23385 12631 23443 12637
rect 23385 12628 23397 12631
rect 20772 12600 23397 12628
rect 20772 12588 20778 12600
rect 23385 12597 23397 12600
rect 23431 12597 23443 12631
rect 23584 12628 23612 12668
rect 25130 12628 25136 12640
rect 23584 12600 25136 12628
rect 23385 12591 23443 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 25406 12588 25412 12640
rect 25464 12588 25470 12640
rect 1104 12538 26220 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 26220 12538
rect 1104 12464 26220 12486
rect 2590 12384 2596 12436
rect 2648 12424 2654 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 2648 12396 3433 12424
rect 2648 12384 2654 12396
rect 3421 12393 3433 12396
rect 3467 12424 3479 12427
rect 5169 12427 5227 12433
rect 3467 12396 5120 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 3602 12316 3608 12368
rect 3660 12356 3666 12368
rect 5092 12356 5120 12396
rect 5169 12393 5181 12427
rect 5215 12424 5227 12427
rect 5626 12424 5632 12436
rect 5215 12396 5632 12424
rect 5215 12393 5227 12396
rect 5169 12387 5227 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 8938 12384 8944 12436
rect 8996 12384 9002 12436
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19668 12396 19901 12424
rect 19668 12384 19674 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 19889 12387 19947 12393
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20533 12427 20591 12433
rect 20533 12424 20545 12427
rect 20220 12396 20545 12424
rect 20220 12384 20226 12396
rect 20533 12393 20545 12396
rect 20579 12393 20591 12427
rect 23566 12424 23572 12436
rect 20533 12387 20591 12393
rect 22204 12396 23572 12424
rect 12897 12359 12955 12365
rect 12897 12356 12909 12359
rect 3660 12328 4016 12356
rect 5092 12328 5672 12356
rect 3660 12316 3666 12328
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 2924 12260 3832 12288
rect 2924 12248 2930 12260
rect 3804 12229 3832 12260
rect 3988 12229 4016 12328
rect 5644 12300 5672 12328
rect 12406 12328 12909 12356
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 9030 12288 9036 12300
rect 7248 12260 9036 12288
rect 7248 12248 7254 12260
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9490 12288 9496 12300
rect 9263 12260 9496 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2363 12192 2789 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 3789 12223 3847 12229
rect 2777 12183 2835 12189
rect 2884 12192 3648 12220
rect 1394 12112 1400 12164
rect 1452 12152 1458 12164
rect 1452 12124 2636 12152
rect 1452 12112 1458 12124
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2133 12087 2191 12093
rect 2133 12084 2145 12087
rect 2004 12056 2145 12084
rect 2004 12044 2010 12056
rect 2133 12053 2145 12056
rect 2179 12053 2191 12087
rect 2133 12047 2191 12053
rect 2406 12044 2412 12096
rect 2464 12044 2470 12096
rect 2498 12044 2504 12096
rect 2556 12044 2562 12096
rect 2608 12084 2636 12124
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 2884 12152 2912 12192
rect 2740 12124 2912 12152
rect 2740 12112 2746 12124
rect 2958 12112 2964 12164
rect 3016 12112 3022 12164
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 3418 12161 3424 12164
rect 3400 12155 3424 12161
rect 3200 12124 3372 12152
rect 3200 12112 3206 12124
rect 3160 12084 3188 12112
rect 2608 12056 3188 12084
rect 3234 12044 3240 12096
rect 3292 12044 3298 12096
rect 3344 12084 3372 12124
rect 3400 12121 3412 12155
rect 3400 12115 3424 12121
rect 3418 12112 3424 12115
rect 3476 12112 3482 12164
rect 3620 12161 3648 12192
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4430 12220 4436 12232
rect 4019 12192 4436 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 5442 12180 5448 12232
rect 5500 12180 5506 12232
rect 8294 12180 8300 12232
rect 8352 12180 8358 12232
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 3605 12155 3663 12161
rect 3605 12121 3617 12155
rect 3651 12152 3663 12155
rect 5169 12155 5227 12161
rect 3651 12124 3832 12152
rect 3651 12121 3663 12124
rect 3605 12115 3663 12121
rect 3804 12096 3832 12124
rect 5169 12121 5181 12155
rect 5215 12152 5227 12155
rect 5258 12152 5264 12164
rect 5215 12124 5264 12152
rect 5215 12121 5227 12124
rect 5169 12115 5227 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 8389 12155 8447 12161
rect 8389 12121 8401 12155
rect 8435 12152 8447 12155
rect 8588 12152 8616 12183
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 9232 12220 9260 12251
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11333 12291 11391 12297
rect 11333 12288 11345 12291
rect 11020 12260 11345 12288
rect 11020 12248 11026 12260
rect 11333 12257 11345 12260
rect 11379 12257 11391 12291
rect 11333 12251 11391 12257
rect 8812 12192 9260 12220
rect 8812 12180 8818 12192
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 11600 12223 11658 12229
rect 11600 12189 11612 12223
rect 11646 12220 11658 12223
rect 12406 12220 12434 12328
rect 12897 12325 12909 12328
rect 12943 12325 12955 12359
rect 20714 12356 20720 12368
rect 12897 12319 12955 12325
rect 20456 12328 20720 12356
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 13136 12260 13461 12288
rect 13136 12248 13142 12260
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 13449 12251 13507 12257
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12257 16267 12291
rect 16209 12251 16267 12257
rect 11646 12192 12434 12220
rect 13265 12223 13323 12229
rect 11646 12189 11658 12192
rect 11600 12183 11658 12189
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13354 12220 13360 12232
rect 13311 12192 13360 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 8435 12124 8616 12152
rect 8435 12121 8447 12124
rect 8389 12115 8447 12121
rect 3694 12084 3700 12096
rect 3344 12056 3700 12084
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 3786 12044 3792 12096
rect 3844 12044 3850 12096
rect 3881 12087 3939 12093
rect 3881 12053 3893 12087
rect 3927 12084 3939 12087
rect 4062 12084 4068 12096
rect 3927 12056 4068 12084
rect 3927 12053 3939 12056
rect 3881 12047 3939 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 5810 12084 5816 12096
rect 5408 12056 5816 12084
rect 5408 12044 5414 12056
rect 5810 12044 5816 12056
rect 5868 12084 5874 12096
rect 6730 12084 6736 12096
rect 5868 12056 6736 12084
rect 5868 12044 5874 12056
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 12713 12087 12771 12093
rect 12713 12053 12725 12087
rect 12759 12084 12771 12087
rect 13280 12084 13308 12183
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 14734 12220 14740 12232
rect 14139 12192 14740 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 16224 12220 16252 12251
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 16908 12260 17877 12288
rect 16908 12248 16914 12260
rect 17865 12257 17877 12260
rect 17911 12288 17923 12291
rect 19794 12288 19800 12300
rect 17911 12260 19800 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 20254 12288 20260 12300
rect 20088 12260 20260 12288
rect 14884 12192 16252 12220
rect 18785 12223 18843 12229
rect 14884 12180 14890 12192
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 14360 12155 14418 12161
rect 14360 12121 14372 12155
rect 14406 12152 14418 12155
rect 14550 12152 14556 12164
rect 14406 12124 14556 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 17681 12155 17739 12161
rect 17681 12121 17693 12155
rect 17727 12152 17739 12155
rect 18141 12155 18199 12161
rect 18141 12152 18153 12155
rect 17727 12124 18153 12152
rect 17727 12121 17739 12124
rect 17681 12115 17739 12121
rect 18141 12121 18153 12124
rect 18187 12121 18199 12155
rect 18141 12115 18199 12121
rect 12759 12056 13308 12084
rect 13357 12087 13415 12093
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 13357 12053 13369 12087
rect 13403 12084 13415 12087
rect 14182 12084 14188 12096
rect 13403 12056 14188 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14516 12056 15485 12084
rect 14516 12044 14522 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15620 12056 15669 12084
rect 15620 12044 15626 12056
rect 15657 12053 15669 12056
rect 15703 12053 15715 12087
rect 15657 12047 15715 12053
rect 16022 12044 16028 12096
rect 16080 12044 16086 12096
rect 16117 12087 16175 12093
rect 16117 12053 16129 12087
rect 16163 12084 16175 12087
rect 16574 12084 16580 12096
rect 16163 12056 16580 12084
rect 16163 12053 16175 12056
rect 16117 12047 16175 12053
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 17310 12044 17316 12096
rect 17368 12044 17374 12096
rect 17770 12044 17776 12096
rect 17828 12044 17834 12096
rect 18800 12084 18828 12183
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 20088 12229 20116 12260
rect 20254 12248 20260 12260
rect 20312 12248 20318 12300
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19760 12192 20085 12220
rect 19760 12180 19766 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20180 12152 20208 12183
rect 20346 12180 20352 12232
rect 20404 12180 20410 12232
rect 20456 12229 20484 12328
rect 20714 12316 20720 12328
rect 20772 12316 20778 12368
rect 21450 12356 21456 12368
rect 20824 12328 21456 12356
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12189 20499 12223
rect 20441 12183 20499 12189
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 20824 12229 20852 12328
rect 21450 12316 21456 12328
rect 21508 12316 21514 12368
rect 22005 12359 22063 12365
rect 22005 12325 22017 12359
rect 22051 12325 22063 12359
rect 22005 12319 22063 12325
rect 22020 12288 22048 12319
rect 21008 12260 22048 12288
rect 21008 12229 21036 12260
rect 20717 12223 20775 12229
rect 20717 12220 20729 12223
rect 20588 12192 20729 12220
rect 20588 12180 20594 12192
rect 20717 12189 20729 12192
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 20993 12223 21051 12229
rect 20993 12189 21005 12223
rect 21039 12189 21051 12223
rect 20993 12183 21051 12189
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21358 12180 21364 12232
rect 21416 12180 21422 12232
rect 21545 12223 21603 12229
rect 21545 12189 21557 12223
rect 21591 12220 21603 12223
rect 21818 12220 21824 12232
rect 21591 12192 21824 12220
rect 21591 12189 21603 12192
rect 21545 12183 21603 12189
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 22204 12229 22232 12396
rect 23566 12384 23572 12396
rect 23624 12424 23630 12436
rect 24762 12424 24768 12436
rect 23624 12396 24768 12424
rect 23624 12384 23630 12396
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 25038 12384 25044 12436
rect 25096 12384 25102 12436
rect 25130 12384 25136 12436
rect 25188 12384 25194 12436
rect 23474 12316 23480 12368
rect 23532 12356 23538 12368
rect 24394 12356 24400 12368
rect 23532 12328 24400 12356
rect 23532 12316 23538 12328
rect 24394 12316 24400 12328
rect 24452 12356 24458 12368
rect 24452 12328 25544 12356
rect 24452 12316 24458 12328
rect 23492 12288 23520 12316
rect 22388 12260 23520 12288
rect 22388 12229 22416 12260
rect 23842 12248 23848 12300
rect 23900 12288 23906 12300
rect 24302 12288 24308 12300
rect 23900 12260 24308 12288
rect 23900 12248 23906 12260
rect 24302 12248 24308 12260
rect 24360 12248 24366 12300
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 24544 12260 24808 12288
rect 24544 12248 24550 12260
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 22373 12223 22431 12229
rect 22373 12189 22385 12223
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 22557 12223 22615 12229
rect 22557 12189 22569 12223
rect 22603 12220 22615 12223
rect 22646 12220 22652 12232
rect 22603 12192 22652 12220
rect 22603 12189 22615 12192
rect 22557 12183 22615 12189
rect 22646 12180 22652 12192
rect 22704 12180 22710 12232
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 23440 12192 24409 12220
rect 23440 12180 23446 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 22281 12155 22339 12161
rect 20180 12124 21312 12152
rect 19334 12084 19340 12096
rect 18800 12056 19340 12084
rect 19334 12044 19340 12056
rect 19392 12084 19398 12096
rect 20162 12084 20168 12096
rect 19392 12056 20168 12084
rect 19392 12044 19398 12056
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20496 12056 21189 12084
rect 20496 12044 20502 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 21284 12084 21312 12124
rect 22281 12121 22293 12155
rect 22327 12121 22339 12155
rect 22281 12115 22339 12121
rect 22094 12084 22100 12096
rect 21284 12056 22100 12084
rect 21177 12047 21235 12053
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 22296 12084 22324 12115
rect 22922 12112 22928 12164
rect 22980 12152 22986 12164
rect 23845 12155 23903 12161
rect 23845 12152 23857 12155
rect 22980 12124 23857 12152
rect 22980 12112 22986 12124
rect 23845 12121 23857 12124
rect 23891 12121 23903 12155
rect 23845 12115 23903 12121
rect 24029 12155 24087 12161
rect 24029 12121 24041 12155
rect 24075 12121 24087 12155
rect 24029 12115 24087 12121
rect 24213 12155 24271 12161
rect 24213 12121 24225 12155
rect 24259 12152 24271 12155
rect 24596 12152 24624 12183
rect 24670 12180 24676 12232
rect 24728 12180 24734 12232
rect 24780 12229 24808 12260
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 24854 12180 24860 12232
rect 24912 12220 24918 12232
rect 25516 12229 25544 12328
rect 25317 12223 25375 12229
rect 25317 12220 25329 12223
rect 24912 12192 25329 12220
rect 24912 12180 24918 12192
rect 25317 12189 25329 12192
rect 25363 12189 25375 12223
rect 25317 12183 25375 12189
rect 25501 12223 25559 12229
rect 25501 12189 25513 12223
rect 25547 12189 25559 12223
rect 25501 12183 25559 12189
rect 25682 12180 25688 12232
rect 25740 12180 25746 12232
rect 24259 12124 24624 12152
rect 24259 12121 24271 12124
rect 24213 12115 24271 12121
rect 23198 12084 23204 12096
rect 22296 12056 23204 12084
rect 23198 12044 23204 12056
rect 23256 12044 23262 12096
rect 24044 12084 24072 12115
rect 25406 12112 25412 12164
rect 25464 12112 25470 12164
rect 25424 12084 25452 12112
rect 25590 12084 25596 12096
rect 24044 12056 25596 12084
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 1104 11994 26220 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 26220 11994
rect 1104 11920 26220 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2406 11880 2412 11892
rect 1627 11852 2412 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2406 11840 2412 11852
rect 2464 11840 2470 11892
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2924 11852 3157 11880
rect 2924 11840 2930 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 3313 11883 3371 11889
rect 3313 11849 3325 11883
rect 3359 11880 3371 11883
rect 3694 11880 3700 11892
rect 3359 11852 3700 11880
rect 3359 11849 3371 11852
rect 3313 11843 3371 11849
rect 3694 11840 3700 11852
rect 3752 11880 3758 11892
rect 3970 11880 3976 11892
rect 3752 11852 3976 11880
rect 3752 11840 3758 11852
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 4798 11880 4804 11892
rect 4387 11852 4804 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 3050 11812 3056 11824
rect 1688 11784 3056 11812
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 1688 11753 1716 11784
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 3513 11815 3571 11821
rect 3513 11812 3525 11815
rect 3476 11784 3525 11812
rect 3476 11772 3482 11784
rect 3513 11781 3525 11784
rect 3559 11812 3571 11815
rect 3559 11784 3832 11812
rect 3559 11781 3571 11784
rect 3513 11775 3571 11781
rect 1946 11753 1952 11756
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1940 11744 1952 11753
rect 1907 11716 1952 11744
rect 1673 11707 1731 11713
rect 1940 11707 1952 11716
rect 1596 11676 1624 11707
rect 1946 11704 1952 11707
rect 2004 11704 2010 11756
rect 3804 11753 3832 11784
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 4356 11812 4384 11843
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5258 11880 5264 11892
rect 5123 11852 5264 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 5718 11840 5724 11892
rect 5776 11840 5782 11892
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 8297 11883 8355 11889
rect 8297 11880 8309 11883
rect 7883 11852 8309 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 8297 11849 8309 11852
rect 8343 11880 8355 11883
rect 8478 11880 8484 11892
rect 8343 11852 8484 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12492 11852 12909 11880
rect 12492 11840 12498 11852
rect 12897 11849 12909 11852
rect 12943 11849 12955 11883
rect 12897 11843 12955 11849
rect 3936 11784 4384 11812
rect 3936 11772 3942 11784
rect 4430 11772 4436 11824
rect 4488 11812 4494 11824
rect 8205 11815 8263 11821
rect 4488 11784 4936 11812
rect 4488 11772 4494 11784
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3804 11676 3832 11707
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 4028 11716 4261 11744
rect 4028 11704 4034 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4706 11744 4712 11756
rect 4571 11716 4712 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4540 11676 4568 11707
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 4908 11753 4936 11784
rect 8205 11781 8217 11815
rect 8251 11812 8263 11815
rect 8754 11812 8760 11824
rect 8251 11784 8760 11812
rect 8251 11781 8263 11784
rect 8205 11775 8263 11781
rect 8754 11772 8760 11784
rect 8812 11772 8818 11824
rect 12912 11812 12940 11843
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 14608 11852 14657 11880
rect 14608 11840 14614 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 19334 11880 19340 11892
rect 18463 11852 19340 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21358 11880 21364 11892
rect 21039 11852 21364 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 25774 11840 25780 11892
rect 25832 11840 25838 11892
rect 12912 11784 13584 11812
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 1596 11648 1716 11676
rect 3804 11648 4568 11676
rect 4617 11679 4675 11685
rect 1688 11540 1716 11648
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 4798 11676 4804 11688
rect 4663 11648 4804 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 3602 11568 3608 11620
rect 3660 11568 3666 11620
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4706 11608 4712 11620
rect 4203 11580 4712 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 4908 11608 4936 11707
rect 5166 11704 5172 11756
rect 5224 11704 5230 11756
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5316 11716 5457 11744
rect 5316 11704 5322 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5552 11676 5580 11707
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 7834 11744 7840 11756
rect 6788 11716 7840 11744
rect 6788 11704 6794 11716
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7892 11716 7941 11744
rect 7892 11704 7898 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8018 11704 8024 11756
rect 8076 11704 8082 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9410 11747 9468 11753
rect 9410 11744 9422 11747
rect 8904 11716 9422 11744
rect 8904 11704 8910 11716
rect 9410 11713 9422 11716
rect 9456 11713 9468 11747
rect 9410 11707 9468 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 10962 11744 10968 11756
rect 9723 11716 10968 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11790 11753 11796 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11020 11716 11529 11744
rect 11020 11704 11026 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11784 11707 11796 11753
rect 11790 11704 11796 11707
rect 11848 11704 11854 11756
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 13188 11753 13216 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13262 11704 13268 11756
rect 13320 11704 13326 11756
rect 5408 11648 5580 11676
rect 5408 11636 5414 11648
rect 7650 11636 7656 11688
rect 7708 11676 7714 11688
rect 8202 11676 8208 11688
rect 7708 11648 8208 11676
rect 7708 11636 7714 11648
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 13004 11676 13032 11704
rect 13004 11648 13216 11676
rect 13188 11620 13216 11648
rect 5261 11611 5319 11617
rect 5261 11608 5273 11611
rect 4908 11580 5273 11608
rect 5261 11577 5273 11580
rect 5307 11577 5319 11611
rect 5261 11571 5319 11577
rect 13170 11568 13176 11620
rect 13228 11568 13234 11620
rect 2958 11540 2964 11552
rect 1688 11512 2964 11540
rect 2958 11500 2964 11512
rect 3016 11540 3022 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 3016 11512 3065 11540
rect 3016 11500 3022 11512
rect 3053 11509 3065 11512
rect 3099 11540 3111 11543
rect 3329 11543 3387 11549
rect 3329 11540 3341 11543
rect 3099 11512 3341 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3329 11509 3341 11512
rect 3375 11540 3387 11543
rect 3878 11540 3884 11552
rect 3375 11512 3884 11540
rect 3375 11509 3387 11512
rect 3329 11503 3387 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 4614 11540 4620 11552
rect 4571 11512 4620 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5626 11540 5632 11552
rect 4856 11512 5632 11540
rect 4856 11500 4862 11512
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 8938 11540 8944 11552
rect 5684 11512 8944 11540
rect 5684 11500 5690 11512
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 13556 11540 13584 11784
rect 13630 11772 13636 11824
rect 13688 11772 13694 11824
rect 17310 11821 17316 11824
rect 17304 11812 17316 11821
rect 14752 11784 17080 11812
rect 17271 11784 17316 11812
rect 14752 11756 14780 11784
rect 17052 11756 17080 11784
rect 17304 11775 17316 11784
rect 17310 11772 17316 11775
rect 17368 11772 17374 11824
rect 20898 11812 20904 11824
rect 19628 11784 20904 11812
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 13964 11716 14289 11744
rect 13964 11704 13970 11716
rect 14277 11713 14289 11716
rect 14323 11744 14335 11747
rect 14458 11744 14464 11756
rect 14323 11716 14464 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14734 11704 14740 11756
rect 14792 11704 14798 11756
rect 15004 11747 15062 11753
rect 15004 11713 15016 11747
rect 15050 11744 15062 11747
rect 15562 11744 15568 11756
rect 15050 11716 15568 11744
rect 15050 11713 15062 11716
rect 15004 11707 15062 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 17034 11704 17040 11756
rect 17092 11704 17098 11756
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19242 11744 19248 11756
rect 18923 11716 19248 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 19628 11753 19656 11784
rect 20898 11772 20904 11784
rect 20956 11812 20962 11824
rect 20956 11784 21864 11812
rect 20956 11772 20962 11784
rect 19886 11753 19892 11756
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 19880 11707 19892 11753
rect 19886 11704 19892 11707
rect 19944 11704 19950 11756
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 21836 11753 21864 11784
rect 23658 11772 23664 11824
rect 23716 11812 23722 11824
rect 24578 11812 24584 11824
rect 23716 11784 24584 11812
rect 23716 11772 23722 11784
rect 24578 11772 24584 11784
rect 24636 11812 24642 11824
rect 24636 11784 24808 11812
rect 24636 11772 24642 11784
rect 21177 11747 21235 11753
rect 21177 11744 21189 11747
rect 20220 11716 21189 11744
rect 20220 11704 20226 11716
rect 21177 11713 21189 11716
rect 21223 11713 21235 11747
rect 21177 11707 21235 11713
rect 21821 11747 21879 11753
rect 21821 11713 21833 11747
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 21910 11704 21916 11756
rect 21968 11744 21974 11756
rect 24118 11753 24124 11756
rect 22077 11747 22135 11753
rect 22077 11744 22089 11747
rect 21968 11716 22089 11744
rect 21968 11704 21974 11716
rect 22077 11713 22089 11716
rect 22123 11713 22135 11747
rect 22077 11707 22135 11713
rect 24112 11707 24124 11753
rect 24118 11704 24124 11707
rect 24176 11704 24182 11756
rect 24780 11744 24808 11784
rect 24780 11716 24900 11744
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 13817 11611 13875 11617
rect 13817 11577 13829 11611
rect 13863 11608 13875 11611
rect 14016 11608 14044 11639
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14240 11648 14780 11676
rect 14240 11636 14246 11648
rect 13863 11580 14044 11608
rect 13863 11577 13875 11580
rect 13817 11571 13875 11577
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 13556 11512 13645 11540
rect 13633 11509 13645 11512
rect 13679 11540 13691 11543
rect 14182 11540 14188 11552
rect 13679 11512 14188 11540
rect 13679 11509 13691 11512
rect 13633 11503 13691 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14752 11540 14780 11648
rect 18966 11636 18972 11688
rect 19024 11636 19030 11688
rect 19058 11636 19064 11688
rect 19116 11636 19122 11688
rect 23842 11636 23848 11688
rect 23900 11636 23906 11688
rect 20714 11568 20720 11620
rect 20772 11608 20778 11620
rect 21818 11608 21824 11620
rect 20772 11580 21824 11608
rect 20772 11568 20778 11580
rect 21818 11568 21824 11580
rect 21876 11568 21882 11620
rect 23658 11608 23664 11620
rect 22756 11580 23664 11608
rect 15654 11540 15660 11552
rect 14752 11512 15660 11540
rect 15654 11500 15660 11512
rect 15712 11540 15718 11552
rect 16022 11540 16028 11552
rect 15712 11512 16028 11540
rect 15712 11500 15718 11512
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16574 11540 16580 11552
rect 16163 11512 16580 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16574 11500 16580 11512
rect 16632 11540 16638 11552
rect 17402 11540 17408 11552
rect 16632 11512 17408 11540
rect 16632 11500 16638 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 18506 11500 18512 11552
rect 18564 11500 18570 11552
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 20588 11512 21281 11540
rect 20588 11500 20594 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21269 11503 21327 11509
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22756 11540 22784 11580
rect 23658 11568 23664 11580
rect 23716 11568 23722 11620
rect 24872 11608 24900 11716
rect 25590 11704 25596 11756
rect 25648 11704 25654 11756
rect 25225 11611 25283 11617
rect 25225 11608 25237 11611
rect 24872 11580 25237 11608
rect 25225 11577 25237 11580
rect 25271 11608 25283 11611
rect 25590 11608 25596 11620
rect 25271 11580 25596 11608
rect 25271 11577 25283 11580
rect 25225 11571 25283 11577
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 22152 11512 22784 11540
rect 22152 11500 22158 11512
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 25314 11540 25320 11552
rect 23256 11512 25320 11540
rect 23256 11500 23262 11512
rect 25314 11500 25320 11512
rect 25372 11500 25378 11552
rect 1104 11450 26220 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 26220 11450
rect 1104 11376 26220 11398
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 4798 11336 4804 11348
rect 4019 11308 4804 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5534 11336 5540 11348
rect 5307 11308 5540 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 6932 11308 7236 11336
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 4080 11172 4353 11200
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 3050 11132 3056 11144
rect 2087 11104 3056 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 2308 11067 2366 11073
rect 2308 11033 2320 11067
rect 2354 11064 2366 11067
rect 3234 11064 3240 11076
rect 2354 11036 3240 11064
rect 2354 11033 2366 11036
rect 2308 11027 2366 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3786 11024 3792 11076
rect 3844 11024 3850 11076
rect 3994 11067 4052 11073
rect 3994 11033 4006 11067
rect 4040 11064 4052 11067
rect 4080 11064 4108 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4706 11200 4712 11212
rect 4341 11163 4399 11169
rect 4448 11172 4712 11200
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 4448 11141 4476 11172
rect 4706 11160 4712 11172
rect 4764 11200 4770 11212
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4764 11172 4997 11200
rect 4764 11160 4770 11172
rect 4985 11169 4997 11172
rect 5031 11200 5043 11203
rect 5031 11172 5488 11200
rect 5031 11169 5043 11172
rect 4985 11163 5043 11169
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 5258 11132 5264 11144
rect 4939 11104 5264 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11101 5411 11135
rect 5460 11132 5488 11172
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 5460 11104 6837 11132
rect 5353 11095 5411 11101
rect 6825 11101 6837 11104
rect 6871 11132 6883 11135
rect 6932 11132 6960 11308
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11237 7159 11271
rect 7101 11231 7159 11237
rect 6871 11104 6960 11132
rect 7116 11132 7144 11231
rect 7208 11200 7236 11308
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7340 11308 7389 11336
rect 7340 11296 7346 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 7834 11296 7840 11348
rect 7892 11296 7898 11348
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 8294 11336 8300 11348
rect 8067 11308 8300 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 8846 11336 8852 11348
rect 8803 11308 8852 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 7561 11271 7619 11277
rect 7561 11237 7573 11271
rect 7607 11268 7619 11271
rect 8478 11268 8484 11280
rect 7607 11240 8484 11268
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8588 11268 8616 11299
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11848 11308 11989 11336
rect 11848 11296 11854 11308
rect 11977 11305 11989 11308
rect 12023 11305 12035 11339
rect 11977 11299 12035 11305
rect 12894 11296 12900 11348
rect 12952 11296 12958 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 14240 11308 14289 11336
rect 14240 11296 14246 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 14277 11299 14335 11305
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 14826 11336 14832 11348
rect 14783 11308 14832 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 8938 11268 8944 11280
rect 8588 11240 8944 11268
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 13078 11268 13084 11280
rect 12406 11240 13084 11268
rect 8018 11200 8024 11212
rect 7208 11172 8024 11200
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8570 11200 8576 11212
rect 8404 11172 8576 11200
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7116 11104 8125 11132
rect 6871 11101 6883 11104
rect 6825 11095 6883 11101
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 4040 11036 4108 11064
rect 4040 11033 4052 11036
rect 3994 11027 4052 11033
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 5368 11064 5396 11095
rect 8202 11092 8208 11144
rect 8260 11092 8266 11144
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 4396 11036 5396 11064
rect 5620 11067 5678 11073
rect 4396 11024 4402 11036
rect 5620 11033 5632 11067
rect 5666 11064 5678 11067
rect 5718 11064 5724 11076
rect 5666 11036 5724 11064
rect 5666 11033 5678 11036
rect 5620 11027 5678 11033
rect 5718 11024 5724 11036
rect 5776 11024 5782 11076
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6788 11036 6929 11064
rect 6788 11024 6794 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 6917 11027 6975 11033
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11033 7159 11067
rect 7101 11027 7159 11033
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 7116 10996 7144 11027
rect 7190 11024 7196 11076
rect 7248 11024 7254 11076
rect 7374 11024 7380 11076
rect 7432 11073 7438 11076
rect 7432 11067 7451 11073
rect 7439 11033 7451 11067
rect 7432 11027 7451 11033
rect 7432 11024 7438 11027
rect 7650 11024 7656 11076
rect 7708 11024 7714 11076
rect 8404 11073 8432 11172
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12406 11132 12434 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 14292 11268 14320 11299
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15004 11339 15062 11345
rect 15004 11305 15016 11339
rect 15050 11305 15062 11339
rect 15004 11299 15062 11305
rect 14918 11268 14924 11280
rect 14292 11240 14924 11268
rect 14918 11228 14924 11240
rect 14976 11268 14982 11280
rect 15019 11268 15047 11299
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18472 11308 18705 11336
rect 18472 11296 18478 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 18693 11299 18751 11305
rect 14976 11240 15047 11268
rect 14976 11228 14982 11240
rect 13262 11200 13268 11212
rect 12636 11172 13268 11200
rect 12636 11144 12664 11172
rect 13262 11160 13268 11172
rect 13320 11200 13326 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 13320 11172 14473 11200
rect 13320 11160 13326 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 12207 11104 12434 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12851 11104 13093 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13170 11092 13176 11144
rect 13228 11092 13234 11144
rect 13630 11132 13636 11144
rect 13280 11104 13636 11132
rect 8662 11073 8668 11076
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11033 8447 11067
rect 8389 11027 8447 11033
rect 8605 11067 8668 11073
rect 8605 11033 8617 11067
rect 8651 11033 8668 11067
rect 8605 11027 8668 11033
rect 8662 11024 8668 11027
rect 8720 11024 8726 11076
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12345 11067 12403 11073
rect 12345 11064 12357 11067
rect 12124 11036 12357 11064
rect 12124 11024 12130 11036
rect 12345 11033 12357 11036
rect 12391 11033 12403 11067
rect 12345 11027 12403 11033
rect 12434 11024 12440 11076
rect 12492 11024 12498 11076
rect 7668 10996 7696 11024
rect 7116 10968 7696 10996
rect 7863 10999 7921 11005
rect 7863 10965 7875 10999
rect 7909 10996 7921 10999
rect 8018 10996 8024 11008
rect 7909 10968 8024 10996
rect 7909 10965 7921 10968
rect 7863 10959 7921 10965
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 12452 10996 12480 11024
rect 13280 10996 13308 11104
rect 13630 11092 13636 11104
rect 13688 11132 13694 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13688 11104 14197 11132
rect 13688 11092 13694 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 14476 11064 14504 11163
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14792 11172 15301 11200
rect 14792 11160 14798 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 17313 11203 17371 11209
rect 17313 11200 17325 11203
rect 17092 11172 17325 11200
rect 17092 11160 17098 11172
rect 17313 11169 17325 11172
rect 17359 11169 17371 11203
rect 18708 11200 18736 11299
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 19886 11296 19892 11348
rect 19944 11336 19950 11348
rect 19981 11339 20039 11345
rect 19981 11336 19993 11339
rect 19944 11308 19993 11336
rect 19944 11296 19950 11308
rect 19981 11305 19993 11308
rect 20027 11305 20039 11339
rect 19981 11299 20039 11305
rect 21729 11339 21787 11345
rect 21729 11305 21741 11339
rect 21775 11336 21787 11339
rect 21910 11336 21916 11348
rect 21775 11308 21916 11336
rect 21775 11305 21787 11308
rect 21729 11299 21787 11305
rect 21910 11296 21916 11308
rect 21968 11296 21974 11348
rect 22922 11296 22928 11348
rect 22980 11336 22986 11348
rect 22980 11308 24992 11336
rect 22980 11296 22986 11308
rect 18966 11228 18972 11280
rect 19024 11268 19030 11280
rect 20717 11271 20775 11277
rect 20717 11268 20729 11271
rect 19024 11240 20024 11268
rect 19024 11228 19030 11240
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 18708 11172 19809 11200
rect 17313 11163 17371 11169
rect 19797 11169 19809 11172
rect 19843 11169 19855 11203
rect 19996 11200 20024 11240
rect 20364 11240 20729 11268
rect 20364 11200 20392 11240
rect 20717 11237 20729 11240
rect 20763 11237 20775 11271
rect 22186 11268 22192 11280
rect 20717 11231 20775 11237
rect 22066 11240 22192 11268
rect 19996 11172 20392 11200
rect 19797 11163 19855 11169
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 21358 11200 21364 11212
rect 20588 11172 20944 11200
rect 20588 11160 20594 11172
rect 17580 11135 17638 11141
rect 17580 11101 17592 11135
rect 17626 11132 17638 11135
rect 18506 11132 18512 11144
rect 17626 11104 18512 11132
rect 17626 11101 17638 11104
rect 17580 11095 17638 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 20254 11092 20260 11144
rect 20312 11092 20318 11144
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 14550 11064 14556 11076
rect 14476 11036 14556 11064
rect 14550 11024 14556 11036
rect 14608 11064 14614 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14608 11036 14841 11064
rect 14608 11024 14614 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 15534 11067 15592 11073
rect 15534 11064 15546 11067
rect 15436 11036 15546 11064
rect 15436 11024 15442 11036
rect 15534 11033 15546 11036
rect 15580 11033 15592 11067
rect 15534 11027 15592 11033
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 20364 11064 20392 11095
rect 20438 11092 20444 11144
rect 20496 11092 20502 11144
rect 20916 11141 20944 11172
rect 21008 11172 21364 11200
rect 21008 11141 21036 11172
rect 21358 11160 21364 11172
rect 21416 11160 21422 11212
rect 22066 11200 22094 11240
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 23566 11228 23572 11280
rect 23624 11268 23630 11280
rect 24857 11271 24915 11277
rect 24857 11268 24869 11271
rect 23624 11240 24869 11268
rect 23624 11228 23630 11240
rect 24857 11237 24869 11240
rect 24903 11237 24915 11271
rect 24857 11231 24915 11237
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 22020 11172 22094 11200
rect 22204 11172 22477 11200
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 20640 11064 20668 11095
rect 21174 11092 21180 11144
rect 21232 11092 21238 11144
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11132 21327 11135
rect 21450 11132 21456 11144
rect 21315 11104 21456 11132
rect 21315 11101 21327 11104
rect 21269 11095 21327 11101
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 22020 11141 22048 11172
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21600 11104 22017 11132
rect 21600 11092 21606 11104
rect 22005 11101 22017 11104
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22204 11141 22232 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 23198 11200 23204 11212
rect 22465 11163 22523 11169
rect 22664 11172 23204 11200
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 22664 11141 22692 11172
rect 23198 11160 23204 11172
rect 23256 11160 23262 11212
rect 23382 11160 23388 11212
rect 23440 11200 23446 11212
rect 23440 11172 23612 11200
rect 23440 11160 23446 11172
rect 23584 11141 23612 11172
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 24213 11203 24271 11209
rect 23716 11172 23888 11200
rect 23716 11160 23722 11172
rect 23860 11141 23888 11172
rect 24213 11169 24225 11203
rect 24259 11169 24271 11203
rect 24964 11200 24992 11308
rect 25774 11296 25780 11348
rect 25832 11296 25838 11348
rect 24213 11163 24271 11169
rect 24780 11172 25268 11200
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11101 23811 11135
rect 23753 11095 23811 11101
rect 23845 11135 23903 11141
rect 23845 11101 23857 11135
rect 23891 11101 23903 11135
rect 23845 11095 23903 11101
rect 21818 11064 21824 11076
rect 17460 11036 20576 11064
rect 20640 11036 21824 11064
rect 17460 11024 17466 11036
rect 12452 10968 13308 10996
rect 14918 10956 14924 11008
rect 14976 10996 14982 11008
rect 15029 10999 15087 11005
rect 15029 10996 15041 10999
rect 14976 10968 15041 10996
rect 14976 10956 14982 10968
rect 15029 10965 15041 10968
rect 15075 10965 15087 10999
rect 15029 10959 15087 10965
rect 15197 10999 15255 11005
rect 15197 10965 15209 10999
rect 15243 10996 15255 10999
rect 15930 10996 15936 11008
rect 15243 10968 15936 10996
rect 15243 10965 15255 10968
rect 15197 10959 15255 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 16669 10999 16727 11005
rect 16669 10965 16681 10999
rect 16715 10996 16727 10999
rect 17126 10996 17132 11008
rect 16715 10968 17132 10996
rect 16715 10965 16727 10968
rect 16669 10959 16727 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 20548 10996 20576 11036
rect 21008 11008 21036 11036
rect 21818 11024 21824 11036
rect 21876 11024 21882 11076
rect 22833 11067 22891 11073
rect 22833 11033 22845 11067
rect 22879 11064 22891 11067
rect 22922 11064 22928 11076
rect 22879 11036 22928 11064
rect 22879 11033 22891 11036
rect 22833 11027 22891 11033
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 23768 11064 23796 11095
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24228 11132 24256 11163
rect 24780 11141 24808 11172
rect 24176 11104 24256 11132
rect 24765 11135 24823 11141
rect 24176 11092 24182 11104
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 23768 11036 24409 11064
rect 24397 11033 24409 11036
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 24578 11024 24584 11076
rect 24636 11024 24642 11076
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 25240 11073 25268 11172
rect 25314 11092 25320 11144
rect 25372 11132 25378 11144
rect 25593 11135 25651 11141
rect 25593 11132 25605 11135
rect 25372 11104 25605 11132
rect 25372 11092 25378 11104
rect 25593 11101 25605 11104
rect 25639 11101 25651 11135
rect 25593 11095 25651 11101
rect 25041 11067 25099 11073
rect 25041 11064 25053 11067
rect 24912 11036 25053 11064
rect 24912 11024 24918 11036
rect 25041 11033 25053 11036
rect 25087 11033 25099 11067
rect 25041 11027 25099 11033
rect 25225 11067 25283 11073
rect 25225 11033 25237 11067
rect 25271 11033 25283 11067
rect 25225 11027 25283 11033
rect 20622 10996 20628 11008
rect 20548 10968 20628 10996
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 20990 10956 20996 11008
rect 21048 10956 21054 11008
rect 1104 10906 26220 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 26220 10906
rect 1104 10832 26220 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3602 10792 3608 10804
rect 2915 10764 3608 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 3786 10752 3792 10804
rect 3844 10792 3850 10804
rect 5445 10795 5503 10801
rect 3844 10764 4535 10792
rect 3844 10752 3850 10764
rect 3050 10684 3056 10736
rect 3108 10724 3114 10736
rect 4338 10724 4344 10736
rect 3108 10696 4344 10724
rect 3108 10684 3114 10696
rect 3993 10659 4051 10665
rect 3993 10625 4005 10659
rect 4039 10656 4051 10659
rect 4154 10656 4160 10668
rect 4039 10628 4160 10656
rect 4039 10625 4051 10628
rect 3993 10619 4051 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 4264 10665 4292 10696
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10625 4307 10659
rect 4507 10656 4535 10764
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 5718 10792 5724 10804
rect 5491 10764 5724 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 7193 10795 7251 10801
rect 7193 10761 7205 10795
rect 7239 10792 7251 10795
rect 7466 10792 7472 10804
rect 7239 10764 7472 10792
rect 7239 10761 7251 10764
rect 7193 10755 7251 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 7650 10792 7656 10804
rect 7607 10764 7656 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 5534 10684 5540 10736
rect 5592 10733 5598 10736
rect 5592 10727 5655 10733
rect 5592 10693 5609 10727
rect 5643 10693 5655 10727
rect 5592 10687 5655 10693
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 7098 10724 7104 10736
rect 5859 10696 7104 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 5592 10684 5598 10687
rect 5828 10656 5856 10687
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 4507 10628 5856 10656
rect 6825 10659 6883 10665
rect 4249 10619 4307 10625
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 7576 10656 7604 10755
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 12342 10792 12348 10804
rect 11655 10764 12348 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12621 10795 12679 10801
rect 12621 10761 12633 10795
rect 12667 10792 12679 10795
rect 13170 10792 13176 10804
rect 12667 10764 13176 10792
rect 12667 10761 12679 10764
rect 12621 10755 12679 10761
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 14918 10792 14924 10804
rect 14415 10764 14924 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 15378 10752 15384 10804
rect 15436 10752 15442 10804
rect 16482 10752 16488 10804
rect 16540 10792 16546 10804
rect 20070 10792 20076 10804
rect 16540 10764 20076 10792
rect 16540 10752 16546 10764
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 21542 10792 21548 10804
rect 21376 10764 21548 10792
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8674 10727 8732 10733
rect 8674 10724 8686 10727
rect 8536 10696 8686 10724
rect 8536 10684 8542 10696
rect 8674 10693 8686 10696
rect 8720 10693 8732 10727
rect 10962 10724 10968 10736
rect 8674 10687 8732 10693
rect 8956 10696 10968 10724
rect 8956 10665 8984 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 14642 10724 14648 10736
rect 11072 10696 14648 10724
rect 6871 10628 7604 10656
rect 8941 10659 8999 10665
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9732 10628 10241 10656
rect 9732 10616 9738 10628
rect 10229 10625 10241 10628
rect 10275 10656 10287 10659
rect 11072 10656 11100 10696
rect 14642 10684 14648 10696
rect 14700 10724 14706 10736
rect 16666 10724 16672 10736
rect 14700 10696 16672 10724
rect 14700 10684 14706 10696
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 21376 10724 21404 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 22278 10792 22284 10804
rect 22020 10764 22284 10792
rect 22020 10733 22048 10764
rect 22278 10752 22284 10764
rect 22336 10792 22342 10804
rect 22646 10792 22652 10804
rect 22336 10764 22652 10792
rect 22336 10752 22342 10764
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 23658 10752 23664 10804
rect 23716 10792 23722 10804
rect 24670 10792 24676 10804
rect 23716 10764 24676 10792
rect 23716 10752 23722 10764
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 25774 10752 25780 10804
rect 25832 10752 25838 10804
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 17144 10696 21404 10724
rect 21468 10696 21833 10724
rect 17144 10668 17172 10696
rect 10275 10628 11100 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11296 10628 11529 10656
rect 11296 10616 11302 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 6730 10548 6736 10600
rect 6788 10548 6794 10600
rect 11716 10520 11744 10619
rect 12084 10588 12112 10619
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 13722 10588 13728 10600
rect 12084 10560 13728 10588
rect 13722 10548 13728 10560
rect 13780 10588 13786 10600
rect 14292 10588 14320 10619
rect 14550 10616 14556 10668
rect 14608 10616 14614 10668
rect 14826 10616 14832 10668
rect 14884 10616 14890 10668
rect 15749 10659 15807 10665
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 17126 10656 17132 10668
rect 15795 10628 17132 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18966 10656 18972 10668
rect 18371 10628 18972 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 21284 10665 21312 10696
rect 21468 10665 21496 10696
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 22005 10727 22063 10733
rect 22005 10693 22017 10727
rect 22051 10693 22063 10727
rect 22005 10687 22063 10693
rect 22189 10727 22247 10733
rect 22189 10693 22201 10727
rect 22235 10724 22247 10727
rect 23290 10724 23296 10736
rect 22235 10696 23296 10724
rect 22235 10693 22247 10696
rect 22189 10687 22247 10693
rect 23290 10684 23296 10696
rect 23348 10684 23354 10736
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21361 10659 21419 10665
rect 21361 10625 21373 10659
rect 21407 10625 21419 10659
rect 21361 10619 21419 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 21683 10628 22094 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 13780 10560 14320 10588
rect 13780 10548 13786 10560
rect 12066 10520 12072 10532
rect 11716 10492 12072 10520
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 12158 10412 12164 10464
rect 12216 10412 12222 10464
rect 14292 10452 14320 10560
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 15841 10591 15899 10597
rect 15841 10588 15853 10591
rect 15712 10560 15853 10588
rect 15712 10548 15718 10560
rect 15841 10557 15853 10560
rect 15887 10557 15899 10591
rect 15841 10551 15899 10557
rect 15930 10548 15936 10600
rect 15988 10548 15994 10600
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 18601 10591 18659 10597
rect 18601 10557 18613 10591
rect 18647 10588 18659 10591
rect 19058 10588 19064 10600
rect 18647 10560 19064 10588
rect 18647 10557 18659 10560
rect 18601 10551 18659 10557
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 21376 10588 21404 10619
rect 21910 10588 21916 10600
rect 21376 10560 21916 10588
rect 21910 10548 21916 10560
rect 21968 10548 21974 10600
rect 22066 10588 22094 10628
rect 22370 10616 22376 10668
rect 22428 10656 22434 10668
rect 23382 10656 23388 10668
rect 22428 10628 23388 10656
rect 22428 10616 22434 10628
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 23566 10616 23572 10668
rect 23624 10616 23630 10668
rect 23676 10665 23704 10752
rect 24029 10727 24087 10733
rect 24029 10693 24041 10727
rect 24075 10724 24087 10727
rect 24366 10727 24424 10733
rect 24366 10724 24378 10727
rect 24075 10696 24378 10724
rect 24075 10693 24087 10696
rect 24029 10687 24087 10693
rect 24366 10693 24378 10696
rect 24412 10693 24424 10727
rect 24366 10687 24424 10693
rect 23661 10659 23719 10665
rect 23661 10625 23673 10659
rect 23707 10625 23719 10659
rect 23661 10619 23719 10625
rect 23750 10616 23756 10668
rect 23808 10656 23814 10668
rect 24210 10656 24216 10668
rect 23808 10628 24216 10656
rect 23808 10616 23814 10628
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25516 10628 25605 10656
rect 22388 10588 22416 10616
rect 24121 10591 24179 10597
rect 24121 10588 24133 10591
rect 22066 10560 22416 10588
rect 23860 10560 24133 10588
rect 23860 10532 23888 10560
rect 24121 10557 24133 10560
rect 24167 10557 24179 10591
rect 24121 10551 24179 10557
rect 19978 10480 19984 10532
rect 20036 10520 20042 10532
rect 20254 10520 20260 10532
rect 20036 10492 20260 10520
rect 20036 10480 20042 10492
rect 20254 10480 20260 10492
rect 20312 10520 20318 10532
rect 23750 10520 23756 10532
rect 20312 10492 23756 10520
rect 20312 10480 20318 10492
rect 23750 10480 23756 10492
rect 23808 10480 23814 10532
rect 23842 10480 23848 10532
rect 23900 10480 23906 10532
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14292 10424 14657 10452
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 15105 10455 15163 10461
rect 15105 10421 15117 10455
rect 15151 10452 15163 10455
rect 16390 10452 16396 10464
rect 15151 10424 16396 10452
rect 15151 10421 15163 10424
rect 15105 10415 15163 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 17957 10455 18015 10461
rect 17957 10452 17969 10455
rect 17920 10424 17969 10452
rect 17920 10412 17926 10424
rect 17957 10421 17969 10424
rect 18003 10421 18015 10455
rect 17957 10415 18015 10421
rect 20990 10412 20996 10464
rect 21048 10412 21054 10464
rect 24854 10412 24860 10464
rect 24912 10452 24918 10464
rect 25516 10461 25544 10628
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 25501 10455 25559 10461
rect 25501 10452 25513 10455
rect 24912 10424 25513 10452
rect 24912 10412 24918 10424
rect 25501 10421 25513 10424
rect 25547 10421 25559 10455
rect 25501 10415 25559 10421
rect 1104 10362 26220 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 26220 10362
rect 1104 10288 26220 10310
rect 12250 10208 12256 10260
rect 12308 10248 12314 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 12308 10220 12725 10248
rect 12308 10208 12314 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 12713 10211 12771 10217
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 14182 10248 14188 10260
rect 13679 10220 14188 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 14550 10208 14556 10260
rect 14608 10248 14614 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14608 10220 14749 10248
rect 14608 10208 14614 10220
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 14737 10211 14795 10217
rect 18966 10208 18972 10260
rect 19024 10208 19030 10260
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 21600 10220 24409 10248
rect 21600 10208 21606 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 24397 10211 24455 10217
rect 25774 10208 25780 10260
rect 25832 10208 25838 10260
rect 11238 10112 11244 10124
rect 9876 10084 11244 10112
rect 3050 10004 3056 10056
rect 3108 10044 3114 10056
rect 3605 10047 3663 10053
rect 3605 10044 3617 10047
rect 3108 10016 3617 10044
rect 3108 10004 3114 10016
rect 3605 10013 3617 10016
rect 3651 10044 3663 10047
rect 3881 10047 3939 10053
rect 3881 10044 3893 10047
rect 3651 10016 3893 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 3881 10013 3893 10016
rect 3927 10013 3939 10047
rect 3881 10007 3939 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 9876 10053 9904 10084
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 14200 10112 14228 10208
rect 15197 10183 15255 10189
rect 15197 10149 15209 10183
rect 15243 10180 15255 10183
rect 15243 10152 15976 10180
rect 15243 10149 15255 10152
rect 15197 10143 15255 10149
rect 15948 10121 15976 10152
rect 22278 10140 22284 10192
rect 22336 10140 22342 10192
rect 15933 10115 15991 10121
rect 14200 10084 14688 10112
rect 9677 10047 9735 10053
rect 4764 10016 6408 10044
rect 4764 10004 4770 10016
rect 6380 9908 6408 10016
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9861 10047 9919 10053
rect 9861 10013 9873 10047
rect 9907 10013 9919 10047
rect 9861 10007 9919 10013
rect 10413 10047 10471 10053
rect 10413 10013 10425 10047
rect 10459 10044 10471 10047
rect 10962 10044 10968 10056
rect 10459 10016 10968 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 9692 9976 9720 10007
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 13354 10004 13360 10056
rect 13412 10004 13418 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13780 10016 14105 10044
rect 13780 10004 13786 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 14550 10044 14556 10056
rect 14323 10016 14556 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 11054 9976 11060 9988
rect 9692 9948 11060 9976
rect 11054 9936 11060 9948
rect 11112 9936 11118 9988
rect 12434 9936 12440 9988
rect 12492 9976 12498 9988
rect 13601 9979 13659 9985
rect 13601 9976 13613 9979
rect 12492 9948 13613 9976
rect 12492 9936 12498 9948
rect 13601 9945 13613 9948
rect 13647 9945 13659 9979
rect 13601 9939 13659 9945
rect 9674 9908 9680 9920
rect 6380 9880 9680 9908
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9769 9911 9827 9917
rect 9769 9877 9781 9911
rect 9815 9908 9827 9911
rect 9950 9908 9956 9920
rect 9815 9880 9956 9908
rect 9815 9877 9827 9880
rect 9769 9871 9827 9877
rect 9950 9868 9956 9880
rect 10008 9868 10014 9920
rect 13446 9868 13452 9920
rect 13504 9868 13510 9920
rect 13740 9908 13768 10004
rect 13817 9979 13875 9985
rect 13817 9945 13829 9979
rect 13863 9976 13875 9979
rect 14292 9976 14320 10007
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14660 10053 14688 10084
rect 15933 10081 15945 10115
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 19794 10072 19800 10124
rect 19852 10072 19858 10124
rect 20898 10072 20904 10124
rect 20956 10072 20962 10124
rect 24762 10112 24768 10124
rect 24596 10084 24768 10112
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 14936 9976 14964 10007
rect 17586 10004 17592 10056
rect 17644 10004 17650 10056
rect 17862 10053 17868 10056
rect 17856 10044 17868 10053
rect 17823 10016 17868 10044
rect 17856 10007 17868 10016
rect 17862 10004 17868 10007
rect 17920 10004 17926 10056
rect 18414 10004 18420 10056
rect 18472 10044 18478 10056
rect 18782 10044 18788 10056
rect 18472 10016 18788 10044
rect 18472 10004 18478 10016
rect 18782 10004 18788 10016
rect 18840 10044 18846 10056
rect 18840 10016 20208 10044
rect 18840 10004 18846 10016
rect 13863 9948 14320 9976
rect 14384 9948 14964 9976
rect 13863 9945 13875 9948
rect 13817 9939 13875 9945
rect 14384 9908 14412 9948
rect 15194 9936 15200 9988
rect 15252 9976 15258 9988
rect 15654 9976 15660 9988
rect 15252 9948 15660 9976
rect 15252 9936 15258 9948
rect 15654 9936 15660 9948
rect 15712 9976 15718 9988
rect 15749 9979 15807 9985
rect 15749 9976 15761 9979
rect 15712 9948 15761 9976
rect 15712 9936 15718 9948
rect 15749 9945 15761 9948
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 17494 9936 17500 9988
rect 17552 9976 17558 9988
rect 19613 9979 19671 9985
rect 17552 9948 19380 9976
rect 17552 9936 17558 9948
rect 13740 9880 14412 9908
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14642 9908 14648 9920
rect 14507 9880 14648 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 15841 9911 15899 9917
rect 15841 9877 15853 9911
rect 15887 9908 15899 9911
rect 16482 9908 16488 9920
rect 15887 9880 16488 9908
rect 15887 9877 15899 9880
rect 15841 9871 15899 9877
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 19242 9868 19248 9920
rect 19300 9868 19306 9920
rect 19352 9908 19380 9948
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 20073 9979 20131 9985
rect 20073 9976 20085 9979
rect 19659 9948 20085 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 20073 9945 20085 9948
rect 20119 9945 20131 9979
rect 20180 9976 20208 10016
rect 20622 10004 20628 10056
rect 20680 10004 20686 10056
rect 20990 10004 20996 10056
rect 21048 10044 21054 10056
rect 21157 10047 21215 10053
rect 21157 10044 21169 10047
rect 21048 10016 21169 10044
rect 21048 10004 21054 10016
rect 21157 10013 21169 10016
rect 21203 10013 21215 10047
rect 21157 10007 21215 10013
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24596 10053 24624 10084
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24084 10016 24593 10044
rect 24084 10004 24090 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 24673 10047 24731 10053
rect 24673 10013 24685 10047
rect 24719 10044 24731 10047
rect 24854 10044 24860 10056
rect 24719 10016 24860 10044
rect 24719 10013 24731 10016
rect 24673 10007 24731 10013
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25130 10044 25136 10056
rect 24995 10016 25136 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25130 10004 25136 10016
rect 25188 10004 25194 10056
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 22462 9976 22468 9988
rect 20180 9948 22468 9976
rect 20073 9939 20131 9945
rect 22462 9936 22468 9948
rect 22520 9976 22526 9988
rect 23934 9976 23940 9988
rect 22520 9948 23940 9976
rect 22520 9936 22526 9948
rect 23934 9936 23940 9948
rect 23992 9936 23998 9988
rect 24394 9936 24400 9988
rect 24452 9976 24458 9988
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 24452 9948 24777 9976
rect 24452 9936 24458 9948
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 19705 9911 19763 9917
rect 19705 9908 19717 9911
rect 19352 9880 19717 9908
rect 19705 9877 19717 9880
rect 19751 9908 19763 9911
rect 21266 9908 21272 9920
rect 19751 9880 21272 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 25240 9908 25268 10007
rect 25590 10004 25596 10056
rect 25648 10004 25654 10056
rect 23532 9880 25268 9908
rect 23532 9868 23538 9880
rect 25406 9868 25412 9920
rect 25464 9868 25470 9920
rect 1104 9818 26220 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 26220 9818
rect 1104 9744 26220 9766
rect 19613 9707 19671 9713
rect 19613 9673 19625 9707
rect 19659 9673 19671 9707
rect 19613 9667 19671 9673
rect 22097 9707 22155 9713
rect 22097 9673 22109 9707
rect 22143 9704 22155 9707
rect 22370 9704 22376 9716
rect 22143 9676 22376 9704
rect 22143 9673 22155 9676
rect 22097 9667 22155 9673
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 3297 9639 3355 9645
rect 3297 9636 3309 9639
rect 1820 9608 3309 9636
rect 1820 9596 1826 9608
rect 3297 9605 3309 9608
rect 3343 9605 3355 9639
rect 3297 9599 3355 9605
rect 3513 9639 3571 9645
rect 3513 9605 3525 9639
rect 3559 9605 3571 9639
rect 11784 9639 11842 9645
rect 3513 9599 3571 9605
rect 9968 9608 11008 9636
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 3528 9500 3556 9599
rect 9968 9577 9996 9608
rect 10980 9580 11008 9608
rect 11784 9605 11796 9639
rect 11830 9636 11842 9639
rect 12158 9636 12164 9648
rect 11830 9608 12164 9636
rect 11830 9605 11842 9608
rect 11784 9599 11842 9605
rect 12158 9596 12164 9608
rect 12216 9596 12222 9648
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 15102 9636 15108 9648
rect 14507 9608 15108 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 15280 9639 15338 9645
rect 15280 9605 15292 9639
rect 15326 9636 15338 9639
rect 15378 9636 15384 9648
rect 15326 9608 15384 9636
rect 15326 9605 15338 9608
rect 15280 9599 15338 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 17856 9639 17914 9645
rect 16448 9608 17264 9636
rect 16448 9596 16454 9608
rect 10226 9577 10232 9580
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9537 10011 9571
rect 10220 9568 10232 9577
rect 10187 9540 10232 9568
rect 9953 9531 10011 9537
rect 10220 9531 10232 9540
rect 2648 9472 3556 9500
rect 2648 9460 2654 9472
rect 2958 9392 2964 9444
rect 3016 9432 3022 9444
rect 4080 9432 4108 9531
rect 10226 9528 10232 9531
rect 10284 9528 10290 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11020 9540 11529 9568
rect 11020 9528 11026 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 14734 9528 14740 9580
rect 14792 9568 14798 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14792 9540 15025 9568
rect 14792 9528 14798 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15120 9568 15148 9596
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 15120 9540 17049 9568
rect 15013 9531 15071 9537
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 9582 9500 9588 9512
rect 9355 9472 9588 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12912 9472 13001 9500
rect 4890 9432 4896 9444
rect 3016 9404 4896 9432
rect 3016 9392 3022 9404
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 12912 9376 12940 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 14642 9460 14648 9512
rect 14700 9460 14706 9512
rect 16482 9500 16488 9512
rect 16408 9472 16488 9500
rect 16408 9441 16436 9472
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 17236 9509 17264 9608
rect 17856 9605 17868 9639
rect 17902 9636 17914 9639
rect 19242 9636 19248 9648
rect 17902 9608 19248 9636
rect 17902 9605 17914 9608
rect 17856 9599 17914 9605
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19628 9636 19656 9667
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 20070 9636 20076 9648
rect 19628 9608 20076 9636
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 19024 9540 19349 9568
rect 19024 9528 19030 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9568 19763 9571
rect 20162 9568 20168 9580
rect 19751 9540 20168 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 21910 9528 21916 9580
rect 21968 9528 21974 9580
rect 22388 9568 22416 9664
rect 23753 9639 23811 9645
rect 23753 9605 23765 9639
rect 23799 9636 23811 9639
rect 24090 9639 24148 9645
rect 24090 9636 24102 9639
rect 23799 9608 24102 9636
rect 23799 9605 23811 9608
rect 23753 9599 23811 9605
rect 24090 9605 24102 9608
rect 24136 9605 24148 9639
rect 24090 9599 24148 9605
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22388 9540 23121 9568
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 23658 9568 23664 9580
rect 23523 9540 23664 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 16393 9435 16451 9441
rect 16393 9401 16405 9435
rect 16439 9401 16451 9435
rect 16393 9395 16451 9401
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 17144 9432 17172 9463
rect 17586 9460 17592 9512
rect 17644 9460 17650 9512
rect 19245 9503 19303 9509
rect 19245 9469 19257 9503
rect 19291 9500 19303 9503
rect 20622 9500 20628 9512
rect 19291 9472 20628 9500
rect 19291 9469 19303 9472
rect 19245 9463 19303 9469
rect 18969 9435 19027 9441
rect 16632 9404 17264 9432
rect 16632 9392 16638 9404
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2832 9336 3157 9364
rect 2832 9324 2838 9336
rect 3145 9333 3157 9336
rect 3191 9333 3203 9367
rect 3145 9327 3203 9333
rect 3326 9324 3332 9376
rect 3384 9324 3390 9376
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4798 9364 4804 9376
rect 3476 9336 4804 9364
rect 3476 9324 3482 9336
rect 4798 9324 4804 9336
rect 4856 9364 4862 9376
rect 6546 9364 6552 9376
rect 4856 9336 6552 9364
rect 4856 9324 4862 9336
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 9861 9367 9919 9373
rect 9861 9333 9873 9367
rect 9907 9364 9919 9367
rect 11054 9364 11060 9376
rect 9907 9336 11060 9364
rect 9907 9333 9919 9336
rect 9861 9327 9919 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 12158 9364 12164 9376
rect 11379 9336 12164 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12894 9324 12900 9376
rect 12952 9324 12958 9376
rect 13633 9367 13691 9373
rect 13633 9333 13645 9367
rect 13679 9364 13691 9367
rect 13722 9364 13728 9376
rect 13679 9336 13728 9364
rect 13679 9333 13691 9336
rect 13633 9327 13691 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14090 9324 14096 9376
rect 14148 9324 14154 9376
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16540 9336 16681 9364
rect 16540 9324 16546 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 17236 9364 17264 9404
rect 18969 9401 18981 9435
rect 19015 9432 19027 9435
rect 19260 9432 19288 9463
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 23400 9500 23428 9531
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 23842 9528 23848 9580
rect 23900 9528 23906 9580
rect 22060 9472 23428 9500
rect 22060 9460 22066 9472
rect 19334 9432 19340 9444
rect 19015 9404 19340 9432
rect 19015 9401 19027 9404
rect 18969 9395 19027 9401
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 17770 9364 17776 9376
rect 17236 9336 17776 9364
rect 16669 9327 16727 9333
rect 17770 9324 17776 9336
rect 17828 9364 17834 9376
rect 19978 9364 19984 9376
rect 17828 9336 19984 9364
rect 17828 9324 17834 9336
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 20806 9364 20812 9376
rect 20496 9336 20812 9364
rect 20496 9324 20502 9336
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 25222 9324 25228 9376
rect 25280 9324 25286 9376
rect 1104 9274 26220 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 26220 9274
rect 1104 9200 26220 9222
rect 1673 9163 1731 9169
rect 1673 9129 1685 9163
rect 1719 9160 1731 9163
rect 1946 9160 1952 9172
rect 1719 9132 1952 9160
rect 1719 9129 1731 9132
rect 1673 9123 1731 9129
rect 1946 9120 1952 9132
rect 2004 9160 2010 9172
rect 3510 9160 3516 9172
rect 2004 9132 3516 9160
rect 2004 9120 2010 9132
rect 2774 8916 2780 8968
rect 2832 8965 2838 8968
rect 2832 8956 2844 8965
rect 2832 8928 2877 8956
rect 2832 8919 2844 8928
rect 2832 8916 2838 8919
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3160 8965 3188 9132
rect 3510 9120 3516 9132
rect 3568 9160 3574 9172
rect 3568 9132 5396 9160
rect 3568 9120 3574 9132
rect 3602 9052 3608 9104
rect 3660 9092 3666 9104
rect 3660 9064 5304 9092
rect 3660 9052 3666 9064
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 3016 8928 3065 8956
rect 3016 8916 3022 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4706 8956 4712 8968
rect 4111 8928 4712 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 3436 8888 3464 8919
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5276 8965 5304 9064
rect 5368 9024 5396 9132
rect 5442 9120 5448 9172
rect 5500 9160 5506 9172
rect 6454 9160 6460 9172
rect 5500 9132 6460 9160
rect 5500 9120 5506 9132
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 9950 9160 9956 9172
rect 8956 9132 9956 9160
rect 5902 9052 5908 9104
rect 5960 9052 5966 9104
rect 5997 9095 6055 9101
rect 5997 9061 6009 9095
rect 6043 9061 6055 9095
rect 5997 9055 6055 9061
rect 5920 9024 5948 9052
rect 5368 8996 5948 9024
rect 6012 9024 6040 9055
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 6641 9095 6699 9101
rect 6641 9092 6653 9095
rect 6236 9064 6653 9092
rect 6236 9052 6242 9064
rect 6641 9061 6653 9064
rect 6687 9061 6699 9095
rect 6641 9055 6699 9061
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7926 9092 7932 9104
rect 7248 9064 7932 9092
rect 7248 9052 7254 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 6546 9024 6552 9036
rect 6012 8996 6552 9024
rect 5368 8965 5396 8996
rect 6546 8984 6552 8996
rect 6604 9024 6610 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6604 8996 6745 9024
rect 6604 8984 6610 8996
rect 6733 8993 6745 8996
rect 6779 9024 6791 9027
rect 6779 8996 6961 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 5776 8928 6408 8956
rect 5776 8916 5782 8928
rect 4614 8888 4620 8900
rect 3436 8860 4620 8888
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 4890 8848 4896 8900
rect 4948 8848 4954 8900
rect 5077 8891 5135 8897
rect 5077 8857 5089 8891
rect 5123 8888 5135 8891
rect 5534 8888 5540 8900
rect 5123 8860 5540 8888
rect 5123 8857 5135 8860
rect 5077 8851 5135 8857
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 5626 8848 5632 8900
rect 5684 8848 5690 8900
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 6273 8891 6331 8897
rect 6273 8888 6285 8891
rect 5960 8860 6285 8888
rect 5960 8848 5966 8860
rect 6273 8857 6285 8860
rect 6319 8857 6331 8891
rect 6380 8888 6408 8928
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6822 8956 6828 8968
rect 6564 8928 6828 8956
rect 6564 8888 6592 8928
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 6933 8965 6961 8996
rect 8956 8965 8984 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 12894 9160 12900 9172
rect 12406 9132 12900 9160
rect 9217 9095 9275 9101
rect 9217 9061 9229 9095
rect 9263 9061 9275 9095
rect 9217 9055 9275 9061
rect 9232 9024 9260 9055
rect 9232 8996 9444 9024
rect 6918 8959 6976 8965
rect 6918 8925 6930 8959
rect 6964 8925 6976 8959
rect 6918 8919 6976 8925
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 6380 8860 6592 8888
rect 9217 8891 9275 8897
rect 6273 8851 6331 8857
rect 9217 8857 9229 8891
rect 9263 8888 9275 8891
rect 9416 8888 9444 8996
rect 12158 8984 12164 9036
rect 12216 8984 12222 9036
rect 12278 9027 12336 9033
rect 12278 8993 12290 9027
rect 12324 9024 12336 9027
rect 12406 9024 12434 9132
rect 12894 9120 12900 9132
rect 12952 9160 12958 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 12952 9132 13277 9160
rect 12952 9120 12958 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 13630 9120 13636 9172
rect 13688 9120 13694 9172
rect 16574 9120 16580 9172
rect 16632 9120 16638 9172
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 19024 9132 19441 9160
rect 19024 9120 19030 9132
rect 19429 9129 19441 9132
rect 19475 9129 19487 9163
rect 22557 9163 22615 9169
rect 22557 9160 22569 9163
rect 19429 9123 19487 9129
rect 20824 9132 22569 9160
rect 12324 8996 12434 9024
rect 13173 9027 13231 9033
rect 12324 8993 12336 8996
rect 12278 8987 12336 8993
rect 13173 8993 13185 9027
rect 13219 9024 13231 9027
rect 13219 8996 14320 9024
rect 13219 8993 13231 8996
rect 13173 8987 13231 8993
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11572 8928 11805 8956
rect 11572 8916 11578 8928
rect 11793 8925 11805 8928
rect 11839 8925 11851 8959
rect 12176 8956 12204 8984
rect 13188 8956 13216 8987
rect 12176 8928 13216 8956
rect 13265 8959 13323 8965
rect 11793 8919 11851 8925
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13630 8956 13636 8968
rect 13495 8928 13636 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 9554 8891 9612 8897
rect 9554 8888 9566 8891
rect 9263 8860 9352 8888
rect 9416 8860 9566 8888
rect 9263 8857 9275 8860
rect 9217 8851 9275 8857
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 3418 8820 3424 8832
rect 3283 8792 3424 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3605 8823 3663 8829
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 4706 8820 4712 8832
rect 3651 8792 4712 8820
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 6181 8823 6239 8829
rect 6181 8820 6193 8823
rect 5776 8792 6193 8820
rect 5776 8780 5782 8792
rect 6181 8789 6193 8792
rect 6227 8820 6239 8823
rect 6730 8820 6736 8832
rect 6227 8792 6736 8820
rect 6227 8789 6239 8792
rect 6181 8783 6239 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 9324 8820 9352 8860
rect 9554 8857 9566 8860
rect 9600 8857 9612 8891
rect 9554 8851 9612 8857
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10781 8891 10839 8897
rect 10781 8888 10793 8891
rect 10560 8860 10793 8888
rect 10560 8848 10566 8860
rect 10781 8857 10793 8860
rect 10827 8857 10839 8891
rect 10781 8851 10839 8857
rect 12069 8891 12127 8897
rect 12069 8857 12081 8891
rect 12115 8888 12127 8891
rect 13280 8888 13308 8919
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14292 8965 14320 8996
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 15197 9027 15255 9033
rect 15197 9024 15209 9027
rect 14792 8996 15209 9024
rect 14792 8984 14798 8996
rect 15197 8993 15209 8996
rect 15243 8993 15255 9027
rect 15197 8987 15255 8993
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 19610 9024 19616 9036
rect 17736 8996 19616 9024
rect 17736 8984 17742 8996
rect 19610 8984 19616 8996
rect 19668 9024 19674 9036
rect 20530 9024 20536 9036
rect 19668 8996 20536 9024
rect 19668 8984 19674 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13872 8928 14105 8956
rect 13872 8916 13878 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 15464 8959 15522 8965
rect 15464 8925 15476 8959
rect 15510 8956 15522 8959
rect 16482 8956 16488 8968
rect 15510 8928 16488 8956
rect 15510 8925 15522 8928
rect 15464 8919 15522 8925
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 18969 8959 19027 8965
rect 18969 8925 18981 8959
rect 19015 8956 19027 8959
rect 19334 8956 19340 8968
rect 19015 8928 19340 8956
rect 19015 8925 19027 8928
rect 18969 8919 19027 8925
rect 19334 8916 19340 8928
rect 19392 8956 19398 8968
rect 19392 8928 19472 8956
rect 19392 8916 19398 8928
rect 13538 8888 13544 8900
rect 12115 8860 12940 8888
rect 13280 8860 13544 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 10226 8820 10232 8832
rect 9324 8792 10232 8820
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 10689 8823 10747 8829
rect 10689 8789 10701 8823
rect 10735 8820 10747 8823
rect 11238 8820 11244 8832
rect 10735 8792 11244 8820
rect 10735 8789 10747 8792
rect 10689 8783 10747 8789
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 12342 8820 12348 8832
rect 11388 8792 12348 8820
rect 11388 8780 11394 8792
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 12526 8780 12532 8832
rect 12584 8780 12590 8832
rect 12912 8820 12940 8860
rect 13538 8848 13544 8860
rect 13596 8888 13602 8900
rect 14185 8891 14243 8897
rect 14185 8888 14197 8891
rect 13596 8860 14197 8888
rect 13596 8848 13602 8860
rect 14185 8857 14197 8860
rect 14231 8857 14243 8891
rect 14185 8851 14243 8857
rect 18690 8848 18696 8900
rect 18748 8888 18754 8900
rect 19444 8897 19472 8928
rect 20438 8916 20444 8968
rect 20496 8956 20502 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20496 8928 20637 8956
rect 20496 8916 20502 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 20714 8916 20720 8968
rect 20772 8916 20778 8968
rect 20824 8965 20852 9132
rect 22557 9129 22569 9132
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 23290 9120 23296 9172
rect 23348 9160 23354 9172
rect 24765 9163 24823 9169
rect 24765 9160 24777 9163
rect 23348 9132 24777 9160
rect 23348 9120 23354 9132
rect 24765 9129 24777 9132
rect 24811 9129 24823 9163
rect 24765 9123 24823 9129
rect 22094 9052 22100 9104
rect 22152 9092 22158 9104
rect 22465 9095 22523 9101
rect 22465 9092 22477 9095
rect 22152 9064 22477 9092
rect 22152 9052 22158 9064
rect 22465 9061 22477 9064
rect 22511 9092 22523 9095
rect 22511 9064 22784 9092
rect 22511 9061 22523 9064
rect 22465 9055 22523 9061
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21085 9027 21143 9033
rect 21085 9024 21097 9027
rect 20956 8996 21097 9024
rect 20956 8984 20962 8996
rect 21085 8993 21097 8996
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 20993 8959 21051 8965
rect 20993 8925 21005 8959
rect 21039 8956 21051 8959
rect 22370 8956 22376 8968
rect 21039 8928 22376 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 22756 8965 22784 9064
rect 22830 9052 22836 9104
rect 22888 9092 22894 9104
rect 24394 9092 24400 9104
rect 22888 9064 24400 9092
rect 22888 9052 22894 9064
rect 24394 9052 24400 9064
rect 24452 9052 24458 9104
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 25222 9024 25228 9036
rect 23440 8996 24339 9024
rect 23440 8984 23446 8996
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8956 22799 8959
rect 23474 8956 23480 8968
rect 22787 8928 23480 8956
rect 22787 8925 22799 8928
rect 22741 8919 22799 8925
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 24311 8956 24339 8996
rect 24596 8996 25228 9024
rect 24596 8965 24624 8996
rect 25222 8984 25228 8996
rect 25280 8984 25286 9036
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 24311 8928 24409 8956
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24688 8928 25268 8956
rect 19245 8891 19303 8897
rect 19245 8888 19257 8891
rect 18748 8860 19257 8888
rect 18748 8848 18754 8860
rect 19245 8857 19257 8860
rect 19291 8857 19303 8891
rect 19245 8851 19303 8857
rect 19429 8891 19487 8897
rect 19429 8857 19441 8891
rect 19475 8857 19487 8891
rect 19429 8851 19487 8857
rect 20349 8891 20407 8897
rect 20349 8857 20361 8891
rect 20395 8888 20407 8891
rect 21330 8891 21388 8897
rect 21330 8888 21342 8891
rect 20395 8860 21342 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 21330 8857 21342 8860
rect 21376 8857 21388 8891
rect 21330 8851 21388 8857
rect 22922 8848 22928 8900
rect 22980 8848 22986 8900
rect 24688 8888 24716 8928
rect 23676 8860 24716 8888
rect 13262 8820 13268 8832
rect 12912 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8820 18935 8823
rect 19058 8820 19064 8832
rect 18923 8792 19064 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19613 8823 19671 8829
rect 19613 8789 19625 8823
rect 19659 8820 19671 8823
rect 21542 8820 21548 8832
rect 19659 8792 21548 8820
rect 19659 8789 19671 8792
rect 19613 8783 19671 8789
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 22940 8820 22968 8848
rect 23676 8820 23704 8860
rect 25038 8848 25044 8900
rect 25096 8848 25102 8900
rect 25240 8897 25268 8928
rect 25590 8916 25596 8968
rect 25648 8916 25654 8968
rect 25225 8891 25283 8897
rect 25225 8857 25237 8891
rect 25271 8888 25283 8891
rect 25314 8888 25320 8900
rect 25271 8860 25320 8888
rect 25271 8857 25283 8860
rect 25225 8851 25283 8857
rect 25314 8848 25320 8860
rect 25372 8848 25378 8900
rect 22940 8792 23704 8820
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 24857 8823 24915 8829
rect 24857 8820 24869 8823
rect 24544 8792 24869 8820
rect 24544 8780 24550 8792
rect 24857 8789 24869 8792
rect 24903 8789 24915 8823
rect 24857 8783 24915 8789
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 1104 8730 26220 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 26220 8730
rect 1104 8656 26220 8678
rect 1762 8576 1768 8628
rect 1820 8576 1826 8628
rect 2590 8576 2596 8628
rect 2648 8576 2654 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 4709 8619 4767 8625
rect 2823 8588 3188 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 1946 8508 1952 8560
rect 2004 8508 2010 8560
rect 2133 8551 2191 8557
rect 2133 8517 2145 8551
rect 2179 8548 2191 8551
rect 3050 8548 3056 8560
rect 2179 8520 3056 8548
rect 2179 8517 2191 8520
rect 2133 8511 2191 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 2958 8480 2964 8492
rect 2884 8452 2964 8480
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2774 8412 2780 8424
rect 2271 8384 2780 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2884 8421 2912 8452
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3160 8489 3188 8588
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 5810 8616 5816 8628
rect 4755 8588 5816 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6178 8576 6184 8628
rect 6236 8576 6242 8628
rect 8754 8616 8760 8628
rect 8128 8588 8760 8616
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3602 8548 3608 8560
rect 3292 8520 3608 8548
rect 3292 8508 3298 8520
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 4522 8508 4528 8560
rect 4580 8508 4586 8560
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5316 8520 6132 8548
rect 5316 8508 5322 8520
rect 3136 8483 3194 8489
rect 3136 8449 3148 8483
rect 3182 8449 3194 8483
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 3136 8443 3194 8449
rect 3896 8452 4353 8480
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 2884 8344 2912 8375
rect 2516 8316 2912 8344
rect 1946 8236 1952 8288
rect 2004 8276 2010 8288
rect 2516 8276 2544 8316
rect 2004 8248 2544 8276
rect 2593 8279 2651 8285
rect 2004 8236 2010 8248
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 3142 8276 3148 8288
rect 2639 8248 3148 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 3786 8276 3792 8288
rect 3292 8248 3792 8276
rect 3292 8236 3298 8248
rect 3786 8236 3792 8248
rect 3844 8276 3850 8288
rect 3896 8276 3924 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5068 8483 5126 8489
rect 5068 8449 5080 8483
rect 5114 8480 5126 8483
rect 5626 8480 5632 8492
rect 5114 8452 5632 8480
rect 5114 8449 5126 8452
rect 5068 8443 5126 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 6104 8344 6132 8520
rect 6196 8480 6224 8576
rect 7374 8508 7380 8560
rect 7432 8548 7438 8560
rect 8128 8557 8156 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9088 8588 11284 8616
rect 9088 8576 9094 8588
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7432 8520 7941 8548
rect 7432 8508 7438 8520
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 8220 8520 8616 8548
rect 8220 8489 8248 8520
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6196 8452 6561 8480
rect 6549 8449 6561 8452
rect 6595 8480 6607 8483
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6595 8452 6929 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8461 8483 8519 8489
rect 8461 8480 8473 8483
rect 8205 8443 8263 8449
rect 8312 8452 8473 8480
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 7116 8344 7144 8443
rect 7852 8412 7880 8443
rect 8018 8412 8024 8424
rect 7852 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8312 8412 8340 8452
rect 8461 8449 8473 8452
rect 8507 8449 8519 8483
rect 8588 8480 8616 8520
rect 9674 8508 9680 8560
rect 9732 8508 9738 8560
rect 11256 8548 11284 8588
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12710 8616 12716 8628
rect 11572 8588 12716 8616
rect 11572 8576 11578 8588
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13814 8616 13820 8628
rect 13740 8588 13820 8616
rect 12066 8548 12072 8560
rect 11256 8520 12072 8548
rect 12066 8508 12072 8520
rect 12124 8548 12130 8560
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12124 8520 13001 8548
rect 12124 8508 12130 8520
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 13740 8548 13768 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 18509 8619 18567 8625
rect 18509 8585 18521 8619
rect 18555 8585 18567 8619
rect 18509 8579 18567 8585
rect 19797 8619 19855 8625
rect 19797 8585 19809 8619
rect 19843 8616 19855 8619
rect 20254 8616 20260 8628
rect 19843 8588 20260 8616
rect 19843 8585 19855 8588
rect 19797 8579 19855 8585
rect 14182 8548 14188 8560
rect 12989 8511 13047 8517
rect 13372 8520 13768 8548
rect 13832 8520 14188 8548
rect 9306 8480 9312 8492
rect 8588 8452 9312 8480
rect 8461 8443 8519 8449
rect 9306 8440 9312 8452
rect 9364 8480 9370 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 9364 8452 11529 8480
rect 9364 8440 9370 8452
rect 10520 8424 10548 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11773 8483 11831 8489
rect 11773 8480 11785 8483
rect 11664 8452 11785 8480
rect 11664 8440 11670 8452
rect 11773 8449 11785 8452
rect 11819 8449 11831 8483
rect 13173 8483 13231 8489
rect 13173 8480 13185 8483
rect 11773 8443 11831 8449
rect 12912 8452 13185 8480
rect 8128 8384 8340 8412
rect 8128 8353 8156 8384
rect 10502 8372 10508 8424
rect 10560 8372 10566 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11238 8412 11244 8424
rect 10827 8384 11244 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 6104 8316 7144 8344
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8313 8171 8347
rect 8113 8307 8171 8313
rect 9582 8304 9588 8356
rect 9640 8304 9646 8356
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10284 8316 11468 8344
rect 10284 8304 10290 8316
rect 3844 8248 3924 8276
rect 4249 8279 4307 8285
rect 3844 8236 3850 8248
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4614 8276 4620 8288
rect 4295 8248 4620 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4614 8236 4620 8248
rect 4672 8276 4678 8288
rect 5442 8276 5448 8288
rect 4672 8248 5448 8276
rect 4672 8236 4678 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 6362 8236 6368 8288
rect 6420 8236 6426 8288
rect 6454 8236 6460 8288
rect 6512 8276 6518 8288
rect 6733 8279 6791 8285
rect 6733 8276 6745 8279
rect 6512 8248 6745 8276
rect 6512 8236 6518 8248
rect 6733 8245 6745 8248
rect 6779 8276 6791 8279
rect 6822 8276 6828 8288
rect 6779 8248 6828 8276
rect 6779 8245 6791 8248
rect 6733 8239 6791 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 7282 8236 7288 8288
rect 7340 8236 7346 8288
rect 11440 8276 11468 8316
rect 11790 8276 11796 8288
rect 11440 8248 11796 8276
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12158 8236 12164 8288
rect 12216 8276 12222 8288
rect 12434 8276 12440 8288
rect 12216 8248 12440 8276
rect 12216 8236 12222 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 12912 8285 12940 8452
rect 13173 8449 13185 8452
rect 13219 8449 13231 8483
rect 13173 8443 13231 8449
rect 13188 8412 13216 8443
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13372 8489 13400 8520
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 13320 8452 13369 8480
rect 13320 8440 13326 8452
rect 13357 8449 13369 8452
rect 13403 8449 13415 8483
rect 13357 8443 13415 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8449 13507 8483
rect 13449 8443 13507 8449
rect 13464 8412 13492 8443
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13832 8489 13860 8520
rect 14182 8508 14188 8520
rect 14240 8548 14246 8560
rect 14734 8548 14740 8560
rect 14240 8520 14740 8548
rect 14240 8508 14246 8520
rect 14734 8508 14740 8520
rect 14792 8548 14798 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 14792 8520 16037 8548
rect 14792 8508 14798 8520
rect 16025 8517 16037 8520
rect 16071 8548 16083 8551
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 16071 8520 17417 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 17405 8517 17417 8520
rect 17451 8548 17463 8551
rect 17586 8548 17592 8560
rect 17451 8520 17592 8548
rect 17451 8517 17463 8520
rect 17405 8511 17463 8517
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 17773 8551 17831 8557
rect 17773 8517 17785 8551
rect 17819 8548 17831 8551
rect 17862 8548 17868 8560
rect 17819 8520 17868 8548
rect 17819 8517 17831 8520
rect 17773 8511 17831 8517
rect 17862 8508 17868 8520
rect 17920 8548 17926 8560
rect 18414 8548 18420 8560
rect 17920 8520 18420 8548
rect 17920 8508 17926 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 14090 8489 14096 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8449 13875 8483
rect 14084 8480 14096 8489
rect 14051 8452 14096 8480
rect 13817 8443 13875 8449
rect 14084 8443 14096 8452
rect 14090 8440 14096 8443
rect 14148 8440 14154 8492
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14608 8452 15240 8480
rect 14608 8440 14614 8452
rect 13630 8412 13636 8424
rect 13188 8384 13636 8412
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13722 8372 13728 8424
rect 13780 8372 13786 8424
rect 15212 8412 15240 8452
rect 16666 8440 16672 8492
rect 16724 8440 16730 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17678 8480 17684 8492
rect 16908 8452 17684 8480
rect 16908 8440 16914 8452
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 18524 8480 18552 8579
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 20990 8616 20996 8628
rect 20772 8588 20996 8616
rect 20772 8576 20778 8588
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 22186 8576 22192 8628
rect 22244 8616 22250 8628
rect 23014 8616 23020 8628
rect 22244 8588 23020 8616
rect 22244 8576 22250 8588
rect 23014 8576 23020 8588
rect 23072 8616 23078 8628
rect 23382 8616 23388 8628
rect 23072 8588 23388 8616
rect 23072 8576 23078 8588
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 23753 8619 23811 8625
rect 23753 8585 23765 8619
rect 23799 8616 23811 8619
rect 23799 8588 23980 8616
rect 23799 8585 23811 8588
rect 23753 8579 23811 8585
rect 18690 8508 18696 8560
rect 18748 8508 18754 8560
rect 20898 8508 20904 8560
rect 20956 8548 20962 8560
rect 22557 8551 22615 8557
rect 22557 8548 22569 8551
rect 20956 8520 22569 8548
rect 20956 8508 20962 8520
rect 22557 8517 22569 8520
rect 22603 8548 22615 8551
rect 23952 8548 23980 8588
rect 24090 8551 24148 8557
rect 24090 8548 24102 8551
rect 22603 8520 23888 8548
rect 23952 8520 24102 8548
rect 22603 8517 22615 8520
rect 22557 8511 22615 8517
rect 23860 8492 23888 8520
rect 24090 8517 24102 8520
rect 24136 8517 24148 8551
rect 25685 8551 25743 8557
rect 25685 8548 25697 8551
rect 24090 8511 24148 8517
rect 24504 8520 25697 8548
rect 19058 8480 19064 8492
rect 18524 8452 19064 8480
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 20303 8452 21312 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 18414 8412 18420 8424
rect 15212 8384 18420 8412
rect 13354 8304 13360 8356
rect 13412 8344 13418 8356
rect 15212 8353 15240 8384
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 18966 8412 18972 8424
rect 18524 8384 18972 8412
rect 15197 8347 15255 8353
rect 13412 8316 13676 8344
rect 13412 8304 13418 8316
rect 13648 8285 13676 8316
rect 15197 8313 15209 8347
rect 15243 8313 15255 8347
rect 15197 8307 15255 8313
rect 17770 8304 17776 8356
rect 17828 8344 17834 8356
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 17828 8316 18337 8344
rect 17828 8304 17834 8316
rect 18325 8313 18337 8316
rect 18371 8313 18383 8347
rect 18325 8307 18383 8313
rect 18524 8285 18552 8384
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 21284 8412 21312 8452
rect 21358 8440 21364 8492
rect 21416 8440 21422 8492
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21600 8452 22017 8480
rect 21600 8440 21606 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 22189 8483 22247 8489
rect 22189 8449 22201 8483
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22204 8412 22232 8443
rect 22370 8440 22376 8492
rect 22428 8440 22434 8492
rect 23106 8440 23112 8492
rect 23164 8440 23170 8492
rect 23293 8483 23351 8489
rect 23293 8449 23305 8483
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 22830 8412 22836 8424
rect 21284 8384 22836 8412
rect 22830 8372 22836 8384
rect 22888 8372 22894 8424
rect 23308 8412 23336 8443
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 23750 8480 23756 8492
rect 23523 8452 23756 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 23750 8440 23756 8452
rect 23808 8440 23814 8492
rect 23842 8440 23848 8492
rect 23900 8440 23906 8492
rect 24504 8480 24532 8520
rect 25685 8517 25697 8520
rect 25731 8517 25743 8551
rect 25685 8511 25743 8517
rect 23952 8452 24532 8480
rect 23952 8412 23980 8452
rect 25314 8440 25320 8492
rect 25372 8440 25378 8492
rect 25501 8483 25559 8489
rect 25501 8449 25513 8483
rect 25547 8480 25559 8483
rect 25590 8480 25596 8492
rect 25547 8452 25596 8480
rect 25547 8449 25559 8452
rect 25501 8443 25559 8449
rect 25516 8412 25544 8443
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 23308 8384 23980 8412
rect 25240 8384 25544 8412
rect 20990 8304 20996 8356
rect 21048 8344 21054 8356
rect 21545 8347 21603 8353
rect 21545 8344 21557 8347
rect 21048 8316 21557 8344
rect 21048 8304 21054 8316
rect 21545 8313 21557 8316
rect 21591 8344 21603 8347
rect 23474 8344 23480 8356
rect 21591 8316 23480 8344
rect 21591 8313 21603 8316
rect 21545 8307 21603 8313
rect 23474 8304 23480 8316
rect 23532 8304 23538 8356
rect 24854 8304 24860 8356
rect 24912 8344 24918 8356
rect 25240 8353 25268 8384
rect 25225 8347 25283 8353
rect 25225 8344 25237 8347
rect 24912 8316 25237 8344
rect 24912 8304 24918 8316
rect 25225 8313 25237 8316
rect 25271 8313 25283 8347
rect 25225 8307 25283 8313
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 12768 8248 12909 8276
rect 12768 8236 12774 8248
rect 12897 8245 12909 8248
rect 12943 8245 12955 8279
rect 12897 8239 12955 8245
rect 13633 8279 13691 8285
rect 13633 8245 13645 8279
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8245 18567 8279
rect 18509 8239 18567 8245
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 21821 8279 21879 8285
rect 21821 8276 21833 8279
rect 20772 8248 21833 8276
rect 20772 8236 20778 8248
rect 21821 8245 21833 8248
rect 21867 8245 21879 8279
rect 21821 8239 21879 8245
rect 1104 8186 26220 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 26220 8186
rect 1104 8112 26220 8134
rect 2409 8075 2467 8081
rect 2409 8041 2421 8075
rect 2455 8072 2467 8075
rect 2774 8072 2780 8084
rect 2455 8044 2780 8072
rect 2455 8041 2467 8044
rect 2409 8035 2467 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 3142 8032 3148 8084
rect 3200 8032 3206 8084
rect 5626 8032 5632 8084
rect 5684 8032 5690 8084
rect 5810 8032 5816 8084
rect 5868 8032 5874 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7653 8075 7711 8081
rect 7653 8072 7665 8075
rect 7432 8044 7665 8072
rect 7432 8032 7438 8044
rect 7653 8041 7665 8044
rect 7699 8041 7711 8075
rect 7653 8035 7711 8041
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 11572 8044 11713 8072
rect 11572 8032 11578 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 11701 8035 11759 8041
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11977 8075 12035 8081
rect 11977 8072 11989 8075
rect 11848 8044 11989 8072
rect 11848 8032 11854 8044
rect 11977 8041 11989 8044
rect 12023 8041 12035 8075
rect 11977 8035 12035 8041
rect 12161 8075 12219 8081
rect 12161 8041 12173 8075
rect 12207 8041 12219 8075
rect 15194 8072 15200 8084
rect 12161 8035 12219 8041
rect 13832 8044 15200 8072
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 8004 3019 8007
rect 3326 8004 3332 8016
rect 3007 7976 3332 8004
rect 3007 7973 3019 7976
rect 2961 7967 3019 7973
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 4172 7976 5488 8004
rect 2884 7908 3648 7936
rect 2884 7877 2912 7908
rect 3620 7880 3648 7908
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2823 7840 2881 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 2409 7803 2467 7809
rect 2409 7769 2421 7803
rect 2455 7800 2467 7803
rect 2590 7800 2596 7812
rect 2455 7772 2596 7800
rect 2455 7769 2467 7772
rect 2409 7763 2467 7769
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 2314 7732 2320 7744
rect 2271 7704 2320 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 2314 7692 2320 7704
rect 2372 7692 2378 7744
rect 3068 7732 3096 7831
rect 3344 7800 3372 7831
rect 3510 7828 3516 7880
rect 3568 7828 3574 7880
rect 3602 7828 3608 7880
rect 3660 7828 3666 7880
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 3988 7800 4016 7831
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4172 7877 4200 7976
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4387 7908 5181 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5460 7936 5488 7976
rect 5534 7964 5540 8016
rect 5592 8004 5598 8016
rect 6086 8004 6092 8016
rect 5592 7976 6092 8004
rect 5592 7964 5598 7976
rect 6086 7964 6092 7976
rect 6144 8004 6150 8016
rect 6181 8007 6239 8013
rect 6181 8004 6193 8007
rect 6144 7976 6193 8004
rect 6144 7964 6150 7976
rect 6181 7973 6193 7976
rect 6227 7973 6239 8007
rect 6181 7967 6239 7973
rect 7469 8007 7527 8013
rect 7469 7973 7481 8007
rect 7515 7973 7527 8007
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 7469 7967 7527 7973
rect 8220 7976 8953 8004
rect 5718 7936 5724 7948
rect 5460 7908 5724 7936
rect 5169 7899 5227 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 7484 7936 7512 7967
rect 8220 7945 8248 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 12176 8004 12204 8035
rect 11112 7976 12204 8004
rect 11112 7964 11118 7976
rect 5868 7908 7512 7936
rect 8021 7939 8079 7945
rect 5868 7896 5874 7908
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 8067 7908 8217 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 10410 7896 10416 7948
rect 10468 7936 10474 7948
rect 10962 7936 10968 7948
rect 10468 7908 10968 7936
rect 10468 7896 10474 7908
rect 10962 7896 10968 7908
rect 11020 7936 11026 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 11020 7908 11161 7936
rect 11020 7896 11026 7908
rect 11149 7905 11161 7908
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12526 7936 12532 7948
rect 11756 7908 12532 7936
rect 11756 7896 11762 7908
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13262 7936 13268 7948
rect 13127 7908 13268 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4764 7840 4813 7868
rect 4764 7828 4770 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7868 5135 7871
rect 5258 7868 5264 7880
rect 5123 7840 5264 7868
rect 5123 7837 5135 7840
rect 5077 7831 5135 7837
rect 4338 7800 4344 7812
rect 3344 7772 3648 7800
rect 3988 7772 4344 7800
rect 3510 7732 3516 7744
rect 3068 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3620 7732 3648 7772
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 5000 7800 5028 7831
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7868 5411 7871
rect 5902 7868 5908 7880
rect 5399 7840 5908 7868
rect 5399 7837 5411 7840
rect 5353 7831 5411 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6696 7840 6741 7868
rect 6696 7828 6702 7840
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7055 7871 7113 7877
rect 7055 7837 7067 7871
rect 7101 7868 7113 7871
rect 7190 7868 7196 7880
rect 7101 7840 7196 7868
rect 7101 7837 7113 7840
rect 7055 7831 7113 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10502 7868 10508 7880
rect 10367 7840 10508 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10873 7871 10931 7877
rect 10873 7837 10885 7871
rect 10919 7837 10931 7871
rect 10873 7831 10931 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 6362 7800 6368 7812
rect 5000 7772 6368 7800
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 6825 7803 6883 7809
rect 6825 7769 6837 7803
rect 6871 7769 6883 7803
rect 9122 7800 9128 7812
rect 6825 7763 6883 7769
rect 7024 7772 9128 7800
rect 4614 7732 4620 7744
rect 3620 7704 4620 7732
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 5534 7692 5540 7744
rect 5592 7692 5598 7744
rect 5810 7692 5816 7744
rect 5868 7692 5874 7744
rect 6840 7732 6868 7763
rect 7024 7732 7052 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 10076 7803 10134 7809
rect 10076 7769 10088 7803
rect 10122 7800 10134 7803
rect 10689 7803 10747 7809
rect 10689 7800 10701 7803
rect 10122 7772 10701 7800
rect 10122 7769 10134 7772
rect 10076 7763 10134 7769
rect 10689 7769 10701 7772
rect 10735 7769 10747 7803
rect 10689 7763 10747 7769
rect 6840 7704 7052 7732
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7193 7735 7251 7741
rect 7193 7732 7205 7735
rect 7156 7704 7205 7732
rect 7156 7692 7162 7704
rect 7193 7701 7205 7704
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8018 7732 8024 7744
rect 7699 7704 8024 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 8754 7692 8760 7744
rect 8812 7732 8818 7744
rect 10888 7732 10916 7831
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11072 7800 11100 7831
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11793 7871 11851 7877
rect 11793 7868 11805 7871
rect 11296 7840 11805 7868
rect 11296 7828 11302 7840
rect 11793 7837 11805 7840
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 12618 7868 12624 7880
rect 11931 7840 12624 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12618 7828 12624 7840
rect 12676 7868 12682 7880
rect 13096 7868 13124 7899
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 13446 7936 13452 7948
rect 13403 7908 13452 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13832 7868 13860 8044
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 17402 8032 17408 8084
rect 17460 8032 17466 8084
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 19300 8044 19349 8072
rect 19300 8032 19306 8044
rect 19337 8041 19349 8044
rect 19383 8072 19395 8075
rect 20898 8072 20904 8084
rect 19383 8044 20904 8072
rect 19383 8041 19395 8044
rect 19337 8035 19395 8041
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 7973 13967 8007
rect 13909 7967 13967 7973
rect 12676 7840 13124 7868
rect 13464 7840 13860 7868
rect 12676 7828 12682 7840
rect 12066 7800 12072 7812
rect 11020 7772 12072 7800
rect 11020 7760 11026 7772
rect 12066 7760 12072 7772
rect 12124 7809 12130 7812
rect 12124 7803 12187 7809
rect 12124 7769 12141 7803
rect 12175 7800 12187 7803
rect 12175 7772 12217 7800
rect 12175 7769 12187 7772
rect 12124 7763 12187 7769
rect 12124 7760 12130 7763
rect 12342 7760 12348 7812
rect 12400 7760 12406 7812
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13464 7809 13492 7840
rect 13449 7803 13507 7809
rect 13449 7800 13461 7803
rect 12584 7772 13461 7800
rect 12584 7760 12590 7772
rect 13449 7769 13461 7772
rect 13495 7769 13507 7803
rect 13924 7800 13952 7967
rect 18046 7964 18052 8016
rect 18104 8004 18110 8016
rect 20622 8004 20628 8016
rect 18104 7976 20628 8004
rect 18104 7964 18110 7976
rect 20622 7964 20628 7976
rect 20680 7964 20686 8016
rect 17034 7896 17040 7948
rect 17092 7936 17098 7948
rect 20070 7936 20076 7948
rect 17092 7908 18920 7936
rect 17092 7896 17098 7908
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14182 7868 14188 7880
rect 14139 7840 14188 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 17862 7868 17868 7880
rect 17543 7840 17868 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 18892 7877 18920 7908
rect 19260 7908 20076 7936
rect 19260 7877 19288 7908
rect 20070 7896 20076 7908
rect 20128 7896 20134 7948
rect 23934 7936 23940 7948
rect 22940 7908 23940 7936
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 18003 7840 18245 7868
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18923 7840 19257 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20806 7868 20812 7880
rect 20763 7840 20812 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 14338 7803 14396 7809
rect 14338 7800 14350 7803
rect 13924 7772 14350 7800
rect 13449 7763 13507 7769
rect 14338 7769 14350 7772
rect 14384 7769 14396 7803
rect 14338 7763 14396 7769
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15620 7772 16129 7800
rect 15620 7760 15626 7772
rect 16117 7769 16129 7772
rect 16163 7769 16175 7803
rect 16117 7763 16175 7769
rect 17681 7803 17739 7809
rect 17681 7769 17693 7803
rect 17727 7800 17739 7803
rect 17972 7800 18000 7831
rect 17727 7772 18000 7800
rect 18325 7803 18383 7809
rect 17727 7769 17739 7772
rect 17681 7763 17739 7769
rect 18325 7769 18337 7803
rect 18371 7800 18383 7803
rect 18800 7800 18828 7831
rect 19536 7800 19564 7831
rect 20806 7828 20812 7840
rect 20864 7868 20870 7880
rect 22940 7877 22968 7908
rect 23934 7896 23940 7908
rect 23992 7936 23998 7948
rect 24397 7939 24455 7945
rect 24397 7936 24409 7939
rect 23992 7908 24409 7936
rect 23992 7896 23998 7908
rect 24397 7905 24409 7908
rect 24443 7905 24455 7939
rect 24397 7899 24455 7905
rect 22925 7871 22983 7877
rect 22925 7868 22937 7871
rect 20864 7840 22937 7868
rect 20864 7828 20870 7840
rect 22925 7837 22937 7840
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23106 7828 23112 7880
rect 23164 7868 23170 7880
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 23164 7840 23213 7868
rect 23164 7828 23170 7840
rect 23201 7837 23213 7840
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 23385 7871 23443 7877
rect 23385 7837 23397 7871
rect 23431 7837 23443 7871
rect 23385 7831 23443 7837
rect 20990 7809 20996 7812
rect 18371 7772 19564 7800
rect 18371 7769 18383 7772
rect 18325 7763 18383 7769
rect 8812 7704 10916 7732
rect 8812 7692 8818 7704
rect 11422 7692 11428 7744
rect 11480 7732 11486 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 11480 7704 11529 7732
rect 11480 7692 11486 7704
rect 11517 7701 11529 7704
rect 11563 7701 11575 7735
rect 11517 7695 11575 7701
rect 12434 7692 12440 7744
rect 12492 7692 12498 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 13587 7704 15485 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 15473 7701 15485 7704
rect 15519 7732 15531 7735
rect 15838 7732 15844 7744
rect 15519 7704 15844 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16574 7692 16580 7744
rect 16632 7732 16638 7744
rect 17696 7732 17724 7763
rect 16632 7704 17724 7732
rect 16632 7692 16638 7704
rect 19058 7692 19064 7744
rect 19116 7692 19122 7744
rect 19536 7732 19564 7772
rect 20984 7763 20996 7809
rect 20990 7760 20996 7763
rect 21048 7760 21054 7812
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 22189 7803 22247 7809
rect 22189 7800 22201 7803
rect 21876 7772 22201 7800
rect 21876 7760 21882 7772
rect 22189 7769 22201 7772
rect 22235 7769 22247 7803
rect 23400 7800 23428 7831
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7868 23627 7871
rect 23750 7868 23756 7880
rect 23615 7840 23756 7868
rect 23615 7837 23627 7840
rect 23569 7831 23627 7837
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 24486 7868 24492 7880
rect 23860 7840 24492 7868
rect 23860 7800 23888 7840
rect 24486 7828 24492 7840
rect 24544 7828 24550 7880
rect 23400 7772 23888 7800
rect 22189 7763 22247 7769
rect 24026 7760 24032 7812
rect 24084 7800 24090 7812
rect 24642 7803 24700 7809
rect 24642 7800 24654 7803
rect 24084 7772 24654 7800
rect 24084 7760 24090 7772
rect 24642 7769 24654 7772
rect 24688 7769 24700 7803
rect 24642 7763 24700 7769
rect 21266 7732 21272 7744
rect 19536 7704 21272 7732
rect 21266 7692 21272 7704
rect 21324 7692 21330 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22370 7732 22376 7744
rect 22152 7704 22376 7732
rect 22152 7692 22158 7704
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 25682 7692 25688 7744
rect 25740 7732 25746 7744
rect 25777 7735 25835 7741
rect 25777 7732 25789 7735
rect 25740 7704 25789 7732
rect 25740 7692 25746 7704
rect 25777 7701 25789 7704
rect 25823 7701 25835 7735
rect 25777 7695 25835 7701
rect 1104 7642 26220 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 26220 7642
rect 1104 7568 26220 7590
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3844 7500 3893 7528
rect 3844 7488 3850 7500
rect 3881 7497 3893 7500
rect 3927 7497 3939 7531
rect 3881 7491 3939 7497
rect 4338 7488 4344 7540
rect 4396 7488 4402 7540
rect 4614 7488 4620 7540
rect 4672 7488 4678 7540
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 6696 7500 7328 7528
rect 6696 7488 6702 7500
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 4033 7463 4091 7469
rect 4033 7460 4045 7463
rect 3660 7432 4045 7460
rect 3660 7420 3666 7432
rect 4033 7429 4045 7432
rect 4079 7429 4091 7463
rect 4033 7423 4091 7429
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7460 4307 7463
rect 4632 7460 4660 7488
rect 4295 7432 4660 7460
rect 4295 7429 4307 7432
rect 4249 7423 4307 7429
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 7300 7460 7328 7500
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11606 7528 11612 7540
rect 10735 7500 11612 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 16574 7528 16580 7540
rect 12207 7500 16580 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 16758 7528 16764 7540
rect 16715 7500 16764 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 20809 7531 20867 7537
rect 19116 7500 20024 7528
rect 19116 7488 19122 7500
rect 8941 7463 8999 7469
rect 8941 7460 8953 7463
rect 5592 7432 6960 7460
rect 7300 7432 7696 7460
rect 5592 7420 5598 7432
rect 2314 7401 2320 7404
rect 2308 7392 2320 7401
rect 2275 7364 2320 7392
rect 2308 7355 2320 7364
rect 2314 7352 2320 7355
rect 2372 7352 2378 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4614 7392 4620 7404
rect 4571 7364 4620 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6932 7392 6960 7432
rect 6990 7395 7048 7401
rect 6990 7392 7002 7395
rect 6932 7364 7002 7392
rect 6825 7355 6883 7361
rect 6990 7361 7002 7364
rect 7036 7361 7048 7395
rect 6990 7355 7048 7361
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 2004 7296 2053 7324
rect 2004 7284 2010 7296
rect 2041 7293 2053 7296
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 4709 7327 4767 7333
rect 4709 7324 4721 7327
rect 3476 7296 4721 7324
rect 3476 7284 3482 7296
rect 4709 7293 4721 7296
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 3292 7160 3433 7188
rect 3292 7148 3298 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3568 7160 4077 7188
rect 3568 7148 3574 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 6840 7188 6868 7355
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7392 7251 7395
rect 7282 7392 7288 7404
rect 7239 7364 7288 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7668 7401 7696 7432
rect 7852 7432 8953 7460
rect 7852 7404 7880 7432
rect 8941 7429 8953 7432
rect 8987 7429 8999 7463
rect 12434 7460 12440 7472
rect 8941 7423 8999 7429
rect 10980 7432 12440 7460
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7423 7364 7481 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7469 7355 7527 7361
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7668 7324 7696 7355
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 7926 7352 7932 7404
rect 7984 7352 7990 7404
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8168 7364 8217 7392
rect 8168 7352 8174 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8536 7364 8677 7392
rect 8536 7352 8542 7364
rect 8665 7361 8677 7364
rect 8711 7361 8723 7395
rect 8665 7355 8723 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 7668 7296 8309 7324
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 7926 7216 7932 7268
rect 7984 7256 7990 7268
rect 8772 7256 8800 7355
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10870 7392 10876 7404
rect 10551 7364 10876 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10980 7401 11008 7432
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 15562 7460 15568 7472
rect 15120 7432 15568 7460
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 12710 7352 12716 7404
rect 12768 7352 12774 7404
rect 15120 7401 15148 7432
rect 15562 7420 15568 7432
rect 15620 7420 15626 7472
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 19613 7463 19671 7469
rect 19613 7460 19625 7463
rect 18748 7432 19288 7460
rect 18748 7420 18754 7432
rect 19260 7404 19288 7432
rect 19352 7432 19625 7460
rect 15378 7401 15384 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 15372 7355 15384 7401
rect 15378 7352 15384 7355
rect 15436 7352 15442 7404
rect 16850 7352 16856 7404
rect 16908 7352 16914 7404
rect 16942 7352 16948 7404
rect 17000 7352 17006 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7361 17279 7395
rect 17221 7355 17279 7361
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7324 11115 7327
rect 11103 7296 11652 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 7984 7228 8800 7256
rect 7984 7216 7990 7228
rect 8478 7188 8484 7200
rect 6840 7160 8484 7188
rect 4065 7151 4123 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 8772 7188 8800 7228
rect 8619 7160 8800 7188
rect 10704 7188 10732 7287
rect 11624 7268 11652 7296
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11940 7296 11989 7324
rect 11940 7284 11946 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 12124 7296 12357 7324
rect 12124 7284 12130 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7324 12679 7327
rect 13446 7324 13452 7336
rect 12667 7296 13452 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 11330 7216 11336 7268
rect 11388 7216 11394 7268
rect 11606 7216 11612 7268
rect 11664 7216 11670 7268
rect 12529 7259 12587 7265
rect 12529 7256 12541 7259
rect 11900 7228 12541 7256
rect 11900 7188 11928 7228
rect 12529 7225 12541 7228
rect 12575 7225 12587 7259
rect 17144 7256 17172 7355
rect 17236 7324 17264 7355
rect 19150 7352 19156 7404
rect 19208 7352 19214 7404
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 19352 7401 19380 7432
rect 19613 7429 19625 7432
rect 19659 7429 19671 7463
rect 19613 7423 19671 7429
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19484 7364 19533 7392
rect 19484 7352 19490 7364
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 19996 7401 20024 7500
rect 20809 7497 20821 7531
rect 20855 7528 20867 7531
rect 20990 7528 20996 7540
rect 20855 7500 20996 7528
rect 20855 7497 20867 7500
rect 20809 7491 20867 7497
rect 20990 7488 20996 7500
rect 21048 7488 21054 7540
rect 22002 7528 22008 7540
rect 21192 7500 22008 7528
rect 20438 7420 20444 7472
rect 20496 7460 20502 7472
rect 20496 7432 21128 7460
rect 20496 7420 20502 7432
rect 20824 7404 20852 7432
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7392 20039 7395
rect 20349 7395 20407 7401
rect 20349 7392 20361 7395
rect 20027 7364 20361 7392
rect 20027 7361 20039 7364
rect 19981 7355 20039 7361
rect 20349 7361 20361 7364
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 17236 7296 20116 7324
rect 19978 7256 19984 7268
rect 17144 7228 19984 7256
rect 12529 7219 12587 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 10704 7160 11928 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 16485 7191 16543 7197
rect 16485 7157 16497 7191
rect 16531 7188 16543 7191
rect 16942 7188 16948 7200
rect 16531 7160 16948 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 18877 7191 18935 7197
rect 18877 7157 18889 7191
rect 18923 7188 18935 7191
rect 19334 7188 19340 7200
rect 18923 7160 19340 7188
rect 18923 7157 18935 7160
rect 18877 7151 18935 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 20088 7188 20116 7296
rect 20364 7256 20392 7355
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 21100 7401 21128 7432
rect 21192 7401 21220 7500
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 24302 7528 24308 7540
rect 23584 7500 24308 7528
rect 21818 7420 21824 7472
rect 21876 7420 21882 7472
rect 23290 7420 23296 7472
rect 23348 7460 23354 7472
rect 23584 7460 23612 7500
rect 24302 7488 24308 7500
rect 24360 7488 24366 7540
rect 25038 7488 25044 7540
rect 25096 7528 25102 7540
rect 25317 7531 25375 7537
rect 25317 7528 25329 7531
rect 25096 7500 25329 7528
rect 25096 7488 25102 7500
rect 25317 7497 25329 7500
rect 25363 7528 25375 7531
rect 25590 7528 25596 7540
rect 25363 7500 25596 7528
rect 25363 7497 25375 7500
rect 25317 7491 25375 7497
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 25777 7531 25835 7537
rect 25777 7497 25789 7531
rect 25823 7528 25835 7531
rect 26142 7528 26148 7540
rect 25823 7500 26148 7528
rect 25823 7497 25835 7500
rect 25777 7491 25835 7497
rect 26142 7488 26148 7500
rect 26200 7488 26206 7540
rect 23348 7432 23612 7460
rect 23348 7420 23354 7432
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 20990 7284 20996 7336
rect 21048 7324 21054 7336
rect 21192 7324 21220 7355
rect 21048 7296 21220 7324
rect 21284 7324 21312 7355
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 21508 7364 23213 7392
rect 21508 7352 21514 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7361 23443 7395
rect 23385 7355 23443 7361
rect 22462 7324 22468 7336
rect 21284 7296 22468 7324
rect 21048 7284 21054 7296
rect 22462 7284 22468 7296
rect 22520 7284 22526 7336
rect 22646 7284 22652 7336
rect 22704 7284 22710 7336
rect 22186 7256 22192 7268
rect 20364 7228 22192 7256
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 23400 7256 23428 7355
rect 23474 7352 23480 7404
rect 23532 7352 23538 7404
rect 23584 7401 23612 7432
rect 23842 7420 23848 7472
rect 23900 7460 23906 7472
rect 24182 7463 24240 7469
rect 24182 7460 24194 7463
rect 23900 7432 24194 7460
rect 23900 7420 23906 7432
rect 24182 7429 24194 7432
rect 24228 7429 24240 7463
rect 24182 7423 24240 7429
rect 23569 7395 23627 7401
rect 23569 7361 23581 7395
rect 23615 7361 23627 7395
rect 23569 7355 23627 7361
rect 23934 7352 23940 7404
rect 23992 7352 23998 7404
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 24728 7364 25605 7392
rect 24728 7352 24734 7364
rect 25593 7361 25605 7364
rect 25639 7392 25651 7395
rect 25682 7392 25688 7404
rect 25639 7364 25688 7392
rect 25639 7361 25651 7364
rect 25593 7355 25651 7361
rect 25682 7352 25688 7364
rect 25740 7352 25746 7404
rect 23845 7327 23903 7333
rect 23845 7293 23857 7327
rect 23891 7324 23903 7327
rect 24044 7324 24072 7352
rect 23891 7296 24072 7324
rect 23891 7293 23903 7296
rect 23845 7287 23903 7293
rect 23474 7256 23480 7268
rect 23400 7228 23480 7256
rect 23474 7216 23480 7228
rect 23532 7216 23538 7268
rect 20622 7188 20628 7200
rect 20088 7160 20628 7188
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 20898 7188 20904 7200
rect 20763 7160 20904 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 1104 7098 26220 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 26220 7098
rect 1104 7024 26220 7046
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7834 6984 7840 6996
rect 7423 6956 7840 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7834 6944 7840 6956
rect 7892 6984 7898 6996
rect 10781 6987 10839 6993
rect 7892 6956 8800 6984
rect 7892 6944 7898 6956
rect 1946 6808 1952 6860
rect 2004 6808 2010 6860
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 3660 6820 4353 6848
rect 3660 6808 3666 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 8772 6848 8800 6956
rect 10781 6953 10793 6987
rect 10827 6984 10839 6987
rect 11422 6984 11428 6996
rect 10827 6956 11428 6984
rect 10827 6953 10839 6956
rect 10781 6947 10839 6953
rect 11422 6944 11428 6956
rect 11480 6984 11486 6996
rect 11974 6984 11980 6996
rect 11480 6956 11980 6984
rect 11480 6944 11486 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 14274 6944 14280 6996
rect 14332 6984 14338 6996
rect 14921 6987 14979 6993
rect 14921 6984 14933 6987
rect 14332 6956 14933 6984
rect 14332 6944 14338 6956
rect 14921 6953 14933 6956
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 16114 6944 16120 6996
rect 16172 6984 16178 6996
rect 19150 6984 19156 6996
rect 16172 6956 19156 6984
rect 16172 6944 16178 6956
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 19426 6984 19432 6996
rect 19260 6956 19432 6984
rect 11054 6916 11060 6928
rect 10888 6888 11060 6916
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8772 6820 8953 6848
rect 4341 6811 4399 6817
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3878 6780 3884 6792
rect 3292 6752 3884 6780
rect 3292 6740 3298 6752
rect 3878 6740 3884 6752
rect 3936 6780 3942 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4614 6780 4620 6792
rect 4212 6752 4620 6780
rect 4212 6740 4218 6752
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 5868 6752 7113 6780
rect 5868 6740 5874 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9631 6752 9689 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10888 6780 10916 6888
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 17957 6919 18015 6925
rect 15028 6888 16988 6916
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11072 6848 11100 6876
rect 11072 6820 11192 6848
rect 10735 6752 10916 6780
rect 11057 6783 11115 6789
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 2216 6715 2274 6721
rect 2216 6681 2228 6715
rect 2262 6712 2274 6715
rect 2314 6712 2320 6724
rect 2262 6684 2320 6712
rect 2262 6681 2274 6684
rect 2216 6675 2274 6681
rect 2314 6672 2320 6684
rect 2372 6672 2378 6724
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3200 6684 3801 6712
rect 3200 6672 3206 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3789 6675 3847 6681
rect 3896 6684 4077 6712
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 3329 6647 3387 6653
rect 3329 6644 3341 6647
rect 2188 6616 3341 6644
rect 2188 6604 2194 6616
rect 3329 6613 3341 6616
rect 3375 6644 3387 6647
rect 3694 6644 3700 6656
rect 3375 6616 3700 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3694 6604 3700 6616
rect 3752 6644 3758 6656
rect 3896 6644 3924 6684
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 8512 6715 8570 6721
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 8846 6712 8852 6724
rect 8558 6684 8852 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 10502 6672 10508 6724
rect 10560 6712 10566 6724
rect 11072 6712 11100 6743
rect 10560 6684 11100 6712
rect 11164 6712 11192 6820
rect 11330 6789 11336 6792
rect 11324 6780 11336 6789
rect 11291 6752 11336 6780
rect 11324 6743 11336 6752
rect 11330 6740 11336 6743
rect 11388 6740 11394 6792
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13872 6752 14105 6780
rect 13872 6740 13878 6752
rect 14093 6749 14105 6752
rect 14139 6780 14151 6783
rect 14642 6780 14648 6792
rect 14139 6752 14648 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14642 6740 14648 6752
rect 14700 6780 14706 6792
rect 15028 6780 15056 6888
rect 16850 6848 16856 6860
rect 15120 6820 16856 6848
rect 15120 6792 15148 6820
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16960 6848 16988 6888
rect 17957 6885 17969 6919
rect 18003 6916 18015 6919
rect 18598 6916 18604 6928
rect 18003 6888 18604 6916
rect 18003 6885 18015 6888
rect 17957 6879 18015 6885
rect 18598 6876 18604 6888
rect 18656 6876 18662 6928
rect 18874 6848 18880 6860
rect 16960 6820 17172 6848
rect 14700 6752 15056 6780
rect 14700 6740 14706 6752
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 15197 6783 15255 6789
rect 15197 6749 15209 6783
rect 15243 6749 15255 6783
rect 15197 6743 15255 6749
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 11882 6712 11888 6724
rect 11164 6684 11888 6712
rect 10560 6672 10566 6684
rect 11882 6672 11888 6684
rect 11940 6672 11946 6724
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 15212 6712 15240 6743
rect 14332 6684 15240 6712
rect 14332 6672 14338 6684
rect 3752 6616 3924 6644
rect 3752 6604 3758 6616
rect 4614 6604 4620 6656
rect 4672 6644 4678 6656
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 4672 6616 7205 6644
rect 4672 6604 4678 6616
rect 7193 6613 7205 6616
rect 7239 6644 7251 6647
rect 7742 6644 7748 6656
rect 7239 6616 7748 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 8168 6616 9781 6644
rect 8168 6604 8174 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11330 6644 11336 6656
rect 11011 6616 11336 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 14461 6647 14519 6653
rect 14461 6613 14473 6647
rect 14507 6644 14519 6647
rect 14550 6644 14556 6656
rect 14507 6616 14556 6644
rect 14507 6613 14519 6616
rect 14461 6607 14519 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15396 6644 15424 6743
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 17144 6789 17172 6820
rect 18423 6820 18880 6848
rect 17129 6783 17187 6789
rect 17129 6749 17141 6783
rect 17175 6780 17187 6783
rect 18046 6780 18052 6792
rect 17175 6752 18052 6780
rect 17175 6749 17187 6752
rect 17129 6743 17187 6749
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18423 6789 18451 6820
rect 18874 6808 18880 6820
rect 18932 6848 18938 6860
rect 19260 6848 19288 6956
rect 19426 6944 19432 6956
rect 19484 6984 19490 6996
rect 19484 6956 20760 6984
rect 19484 6944 19490 6956
rect 18932 6820 19288 6848
rect 20732 6848 20760 6956
rect 21542 6944 21548 6996
rect 21600 6944 21606 6996
rect 24210 6984 24216 6996
rect 22388 6956 24216 6984
rect 21450 6848 21456 6860
rect 20732 6820 21456 6848
rect 18932 6808 18938 6820
rect 18405 6783 18463 6789
rect 18405 6749 18417 6783
rect 18451 6749 18463 6783
rect 18405 6743 18463 6749
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 18690 6740 18696 6792
rect 18748 6740 18754 6792
rect 18782 6740 18788 6792
rect 18840 6740 18846 6792
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 20732 6789 20760 6820
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 21560 6848 21588 6944
rect 22388 6848 22416 6956
rect 24210 6944 24216 6956
rect 24268 6984 24274 6996
rect 24578 6984 24584 6996
rect 24268 6956 24584 6984
rect 24268 6944 24274 6956
rect 24578 6944 24584 6956
rect 24636 6944 24642 6996
rect 24670 6916 24676 6928
rect 23676 6888 24676 6916
rect 21560 6820 22416 6848
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19208 6752 19257 6780
rect 19208 6740 19214 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 20717 6783 20775 6789
rect 20717 6749 20729 6783
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 20990 6740 20996 6792
rect 21048 6740 21054 6792
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 15562 6672 15568 6724
rect 15620 6712 15626 6724
rect 15841 6715 15899 6721
rect 15841 6712 15853 6715
rect 15620 6684 15853 6712
rect 15620 6672 15626 6684
rect 15841 6681 15853 6684
rect 15887 6681 15899 6715
rect 15841 6675 15899 6681
rect 16850 6672 16856 6724
rect 16908 6712 16914 6724
rect 16945 6715 17003 6721
rect 16945 6712 16957 6715
rect 16908 6684 16957 6712
rect 16908 6672 16914 6684
rect 16945 6681 16957 6684
rect 16991 6681 17003 6715
rect 16945 6675 17003 6681
rect 18141 6715 18199 6721
rect 18141 6681 18153 6715
rect 18187 6681 18199 6715
rect 18141 6675 18199 6681
rect 18325 6715 18383 6721
rect 18325 6681 18337 6715
rect 18371 6712 18383 6715
rect 18966 6712 18972 6724
rect 18371 6684 18972 6712
rect 18371 6681 18383 6684
rect 18325 6675 18383 6681
rect 15930 6644 15936 6656
rect 15396 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16022 6604 16028 6656
rect 16080 6644 16086 6656
rect 16761 6647 16819 6653
rect 16761 6644 16773 6647
rect 16080 6616 16773 6644
rect 16080 6604 16086 6616
rect 16761 6613 16773 6616
rect 16807 6613 16819 6647
rect 16761 6607 16819 6613
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18156 6644 18184 6675
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19061 6715 19119 6721
rect 19061 6681 19073 6715
rect 19107 6712 19119 6715
rect 19490 6715 19548 6721
rect 19490 6712 19502 6715
rect 19107 6684 19502 6712
rect 19107 6681 19119 6684
rect 19061 6675 19119 6681
rect 19490 6681 19502 6684
rect 19536 6681 19548 6715
rect 21100 6712 21128 6743
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 22388 6789 22416 6820
rect 22462 6808 22468 6860
rect 22520 6848 22526 6860
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 22520 6820 22661 6848
rect 22520 6808 22526 6820
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 23474 6808 23480 6860
rect 23532 6808 23538 6860
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21324 6752 22201 6780
rect 21324 6740 21330 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 22922 6780 22928 6792
rect 22603 6752 22928 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 22922 6740 22928 6752
rect 22980 6780 22986 6792
rect 23676 6789 23704 6888
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 23661 6783 23719 6789
rect 22980 6752 23612 6780
rect 22980 6740 22986 6752
rect 21726 6712 21732 6724
rect 21100 6684 21732 6712
rect 19490 6675 19548 6681
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 22833 6715 22891 6721
rect 22833 6712 22845 6715
rect 22152 6684 22845 6712
rect 22152 6672 22158 6684
rect 22833 6681 22845 6684
rect 22879 6681 22891 6715
rect 22833 6675 22891 6681
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 18012 6616 20637 6644
rect 18012 6604 18018 6616
rect 20625 6613 20637 6616
rect 20671 6644 20683 6647
rect 20714 6644 20720 6656
rect 20671 6616 20720 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 21358 6604 21364 6656
rect 21416 6604 21422 6656
rect 22848 6644 22876 6675
rect 23014 6672 23020 6724
rect 23072 6672 23078 6724
rect 23584 6712 23612 6752
rect 23661 6749 23673 6783
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 24578 6740 24584 6792
rect 24636 6740 24642 6792
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 24946 6740 24952 6792
rect 25004 6740 25010 6792
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 23845 6715 23903 6721
rect 23845 6712 23857 6715
rect 23584 6684 23857 6712
rect 23845 6681 23857 6684
rect 23891 6681 23903 6715
rect 23845 6675 23903 6681
rect 23952 6684 24532 6712
rect 23952 6644 23980 6684
rect 22848 6616 23980 6644
rect 24394 6604 24400 6656
rect 24452 6604 24458 6656
rect 24504 6644 24532 6684
rect 24762 6672 24768 6724
rect 24820 6672 24826 6724
rect 25240 6644 25268 6743
rect 25590 6740 25596 6792
rect 25648 6740 25654 6792
rect 24504 6616 25268 6644
rect 25406 6604 25412 6656
rect 25464 6604 25470 6656
rect 25774 6604 25780 6656
rect 25832 6604 25838 6656
rect 1104 6554 26220 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 26220 6554
rect 1104 6480 26220 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6409 2283 6443
rect 2225 6403 2283 6409
rect 2130 6332 2136 6384
rect 2188 6332 2194 6384
rect 2240 6372 2268 6403
rect 2314 6400 2320 6452
rect 2372 6400 2378 6452
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 3881 6443 3939 6449
rect 3881 6440 3893 6443
rect 2976 6412 3893 6440
rect 2469 6375 2527 6381
rect 2469 6372 2481 6375
rect 2240 6344 2481 6372
rect 2469 6341 2481 6344
rect 2515 6341 2527 6375
rect 2469 6335 2527 6341
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 2976 6372 3004 6412
rect 3881 6409 3893 6412
rect 3927 6440 3939 6443
rect 4062 6440 4068 6452
rect 3927 6412 4068 6440
rect 3927 6409 3939 6412
rect 3881 6403 3939 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6454 6440 6460 6452
rect 6043 6412 6460 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6546 6400 6552 6452
rect 6604 6400 6610 6452
rect 8110 6400 8116 6452
rect 8168 6400 8174 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 8941 6443 8999 6449
rect 8941 6440 8953 6443
rect 8904 6412 8953 6440
rect 8904 6400 8910 6412
rect 8941 6409 8953 6412
rect 8987 6409 8999 6443
rect 10962 6440 10968 6452
rect 8941 6403 8999 6409
rect 10888 6412 10968 6440
rect 2731 6344 3004 6372
rect 3068 6344 3740 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 2590 6304 2596 6316
rect 2271 6276 2596 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 1964 6236 1992 6267
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 3068 6313 3096 6344
rect 3712 6316 3740 6344
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 5169 6375 5227 6381
rect 5169 6372 5181 6375
rect 4672 6344 5181 6372
rect 4672 6332 4678 6344
rect 5169 6341 5181 6344
rect 5215 6341 5227 6375
rect 5169 6335 5227 6341
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 5369 6375 5427 6381
rect 5369 6372 5381 6375
rect 5316 6344 5381 6372
rect 5316 6332 5322 6344
rect 5369 6341 5381 6344
rect 5415 6341 5427 6375
rect 6564 6372 6592 6400
rect 7926 6372 7932 6384
rect 5369 6335 5427 6341
rect 5828 6344 6592 6372
rect 7392 6344 7932 6372
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 3234 6264 3240 6316
rect 3292 6264 3298 6316
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 1964 6208 2973 6236
rect 2608 6112 2636 6208
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 3160 6236 3188 6264
rect 3528 6236 3556 6267
rect 3694 6264 3700 6316
rect 3752 6264 3758 6316
rect 5828 6313 5856 6344
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6086 6264 6092 6316
rect 6144 6264 6150 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6454 6304 6460 6316
rect 6411 6276 6460 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 7392 6313 7420 6344
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 9033 6375 9091 6381
rect 9033 6372 9045 6375
rect 8352 6344 9045 6372
rect 8352 6332 8358 6344
rect 9033 6341 9045 6344
rect 9079 6341 9091 6375
rect 9033 6335 9091 6341
rect 9401 6375 9459 6381
rect 9401 6341 9413 6375
rect 9447 6372 9459 6375
rect 9645 6375 9703 6381
rect 9645 6372 9657 6375
rect 9447 6344 9657 6372
rect 9447 6341 9459 6344
rect 9401 6335 9459 6341
rect 9645 6341 9657 6344
rect 9691 6341 9703 6375
rect 9645 6335 9703 6341
rect 9861 6375 9919 6381
rect 9861 6341 9873 6375
rect 9907 6341 9919 6375
rect 9861 6335 9919 6341
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 3160 6208 3556 6236
rect 6104 6236 6132 6264
rect 6564 6236 6592 6267
rect 7466 6264 7472 6316
rect 7524 6264 7530 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8386 6304 8392 6316
rect 8251 6276 8392 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8938 6304 8944 6316
rect 8536 6276 8944 6304
rect 8536 6264 8542 6276
rect 8938 6264 8944 6276
rect 8996 6304 9002 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8996 6276 9229 6304
rect 8996 6264 9002 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9876 6304 9904 6335
rect 10888 6313 10916 6412
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 14182 6440 14188 6452
rect 11020 6412 14188 6440
rect 11020 6400 11026 6412
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15436 6412 15577 6440
rect 15436 6400 15442 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 15988 6412 16681 6440
rect 15988 6400 15994 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 24394 6440 24400 6452
rect 16669 6403 16727 6409
rect 18800 6412 24400 6440
rect 11057 6375 11115 6381
rect 11057 6341 11069 6375
rect 11103 6372 11115 6375
rect 12066 6372 12072 6384
rect 11103 6344 12072 6372
rect 11103 6341 11115 6344
rect 11057 6335 11115 6341
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 13280 6344 14228 6372
rect 9364 6276 9904 6304
rect 10873 6307 10931 6313
rect 9364 6264 9370 6276
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 13280 6313 13308 6344
rect 11195 6307 11253 6313
rect 11195 6273 11207 6307
rect 11241 6304 11253 6307
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11241 6276 11805 6304
rect 11241 6273 11253 6276
rect 11195 6267 11253 6273
rect 11793 6273 11805 6276
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13532 6307 13590 6313
rect 13532 6273 13544 6307
rect 13578 6304 13590 6307
rect 14090 6304 14096 6316
rect 13578 6276 14096 6304
rect 13578 6273 13590 6276
rect 13532 6267 13590 6273
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 14200 6304 14228 6344
rect 15470 6332 15476 6384
rect 15528 6372 15534 6384
rect 18800 6372 18828 6412
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 19334 6381 19340 6384
rect 19328 6372 19340 6381
rect 15528 6344 18828 6372
rect 19295 6344 19340 6372
rect 15528 6332 15534 6344
rect 19328 6335 19340 6344
rect 19334 6332 19340 6335
rect 19392 6332 19398 6384
rect 23569 6375 23627 6381
rect 22066 6344 23428 6372
rect 15562 6304 15568 6316
rect 14200 6276 15568 6304
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 15930 6264 15936 6316
rect 15988 6264 15994 6316
rect 16022 6264 16028 6316
rect 16080 6264 16086 6316
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 6104 6208 6592 6236
rect 7929 6239 7987 6245
rect 2961 6199 3019 6205
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 7975 6208 8309 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 2976 6168 3004 6199
rect 11330 6196 11336 6248
rect 11388 6196 11394 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 12032 6208 12357 6236
rect 12032 6196 12038 6208
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 16224 6236 16252 6267
rect 16758 6264 16764 6316
rect 16816 6304 16822 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16816 6276 16865 6304
rect 16816 6264 16822 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 16942 6264 16948 6316
rect 17000 6264 17006 6316
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 19794 6304 19800 6316
rect 17267 6276 19800 6304
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 21266 6264 21272 6316
rect 21324 6264 21330 6316
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 16390 6236 16396 6248
rect 14792 6208 16396 6236
rect 14792 6196 14798 6208
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 17052 6236 17080 6264
rect 16960 6208 17080 6236
rect 3418 6168 3424 6180
rect 2976 6140 3424 6168
rect 3418 6128 3424 6140
rect 3476 6168 3482 6180
rect 4154 6168 4160 6180
rect 3476 6140 4160 6168
rect 3476 6128 3482 6140
rect 4154 6128 4160 6140
rect 4212 6128 4218 6180
rect 6457 6171 6515 6177
rect 6457 6168 6469 6171
rect 5368 6140 6469 6168
rect 2498 6060 2504 6112
rect 2556 6060 2562 6112
rect 2590 6060 2596 6112
rect 2648 6060 2654 6112
rect 5368 6109 5396 6140
rect 6457 6137 6469 6140
rect 6503 6137 6515 6171
rect 6457 6131 6515 6137
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 8444 6140 9720 6168
rect 8444 6128 8450 6140
rect 5353 6103 5411 6109
rect 5353 6069 5365 6103
rect 5399 6069 5411 6103
rect 5353 6063 5411 6069
rect 5534 6060 5540 6112
rect 5592 6060 5598 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5718 6100 5724 6112
rect 5675 6072 5724 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 7653 6103 7711 6109
rect 7653 6069 7665 6103
rect 7699 6100 7711 6103
rect 8294 6100 8300 6112
rect 7699 6072 8300 6100
rect 7699 6069 7711 6072
rect 7653 6063 7711 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 9692 6109 9720 6140
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 14516 6140 15976 6168
rect 14516 6128 14522 6140
rect 15948 6112 15976 6140
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 16960 6168 16988 6208
rect 19058 6196 19064 6248
rect 19116 6196 19122 6248
rect 20254 6196 20260 6248
rect 20312 6236 20318 6248
rect 21376 6236 21404 6267
rect 21450 6264 21456 6316
rect 21508 6304 21514 6316
rect 21726 6304 21732 6316
rect 21508 6276 21732 6304
rect 21508 6264 21514 6276
rect 21726 6264 21732 6276
rect 21784 6304 21790 6316
rect 22066 6304 22094 6344
rect 21784 6276 22094 6304
rect 22925 6307 22983 6313
rect 21784 6264 21790 6276
rect 22925 6273 22937 6307
rect 22971 6304 22983 6307
rect 23014 6304 23020 6316
rect 22971 6276 23020 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 23106 6264 23112 6316
rect 23164 6264 23170 6316
rect 23198 6264 23204 6316
rect 23256 6264 23262 6316
rect 23290 6264 23296 6316
rect 23348 6264 23354 6316
rect 23400 6304 23428 6344
rect 23569 6341 23581 6375
rect 23615 6372 23627 6375
rect 23906 6375 23964 6381
rect 23906 6372 23918 6375
rect 23615 6344 23918 6372
rect 23615 6341 23627 6344
rect 23569 6335 23627 6341
rect 23906 6341 23918 6344
rect 23952 6341 23964 6375
rect 23906 6335 23964 6341
rect 25409 6375 25467 6381
rect 25409 6341 25421 6375
rect 25455 6372 25467 6375
rect 25590 6372 25596 6384
rect 25455 6344 25596 6372
rect 25455 6341 25467 6344
rect 25409 6335 25467 6341
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 23750 6304 23756 6316
rect 23400 6276 23756 6304
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 24670 6264 24676 6316
rect 24728 6304 24734 6316
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 24728 6276 25329 6304
rect 24728 6264 24734 6276
rect 25317 6273 25329 6276
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 25501 6307 25559 6313
rect 25501 6273 25513 6307
rect 25547 6273 25559 6307
rect 25501 6267 25559 6273
rect 25685 6307 25743 6313
rect 25685 6273 25697 6307
rect 25731 6273 25743 6307
rect 25685 6267 25743 6273
rect 22554 6236 22560 6248
rect 20312 6208 22560 6236
rect 20312 6196 20318 6208
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 22646 6196 22652 6248
rect 22704 6236 22710 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 22704 6208 23673 6236
rect 22704 6196 22710 6208
rect 23661 6205 23673 6208
rect 23707 6205 23719 6239
rect 23661 6199 23719 6205
rect 24762 6196 24768 6248
rect 24820 6236 24826 6248
rect 25516 6236 25544 6267
rect 24820 6208 25544 6236
rect 24820 6196 24826 6208
rect 16264 6140 16988 6168
rect 16264 6128 16270 6140
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 21726 6168 21732 6180
rect 20588 6140 21732 6168
rect 20588 6128 20594 6140
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 24946 6128 24952 6180
rect 25004 6168 25010 6180
rect 25004 6140 25268 6168
rect 25004 6128 25010 6140
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 10778 6100 10784 6112
rect 10735 6072 10784 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14274 6100 14280 6112
rect 13964 6072 14280 6100
rect 13964 6060 13970 6072
rect 14274 6060 14280 6072
rect 14332 6100 14338 6112
rect 14645 6103 14703 6109
rect 14645 6100 14657 6103
rect 14332 6072 14657 6100
rect 14332 6060 14338 6072
rect 14645 6069 14657 6072
rect 14691 6069 14703 6103
rect 14645 6063 14703 6069
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 17402 6100 17408 6112
rect 15988 6072 17408 6100
rect 15988 6060 15994 6072
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20441 6103 20499 6109
rect 20441 6100 20453 6103
rect 19852 6072 20453 6100
rect 19852 6060 19858 6072
rect 20441 6069 20453 6072
rect 20487 6100 20499 6103
rect 20898 6100 20904 6112
rect 20487 6072 20904 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 21542 6060 21548 6112
rect 21600 6060 21606 6112
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 25056 6109 25084 6140
rect 25041 6103 25099 6109
rect 25041 6100 25053 6103
rect 24084 6072 25053 6100
rect 24084 6060 24090 6072
rect 25041 6069 25053 6072
rect 25087 6069 25099 6103
rect 25041 6063 25099 6069
rect 25130 6060 25136 6112
rect 25188 6060 25194 6112
rect 25240 6100 25268 6140
rect 25314 6128 25320 6180
rect 25372 6168 25378 6180
rect 25700 6168 25728 6267
rect 25372 6140 25728 6168
rect 25372 6128 25378 6140
rect 25590 6100 25596 6112
rect 25240 6072 25596 6100
rect 25590 6060 25596 6072
rect 25648 6060 25654 6112
rect 1104 6010 26220 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 26220 6010
rect 1104 5936 26220 5958
rect 2498 5856 2504 5908
rect 2556 5896 2562 5908
rect 4430 5896 4436 5908
rect 2556 5868 4436 5896
rect 2556 5856 2562 5868
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 5258 5896 5264 5908
rect 4847 5868 5264 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 6776 5896
rect 5592 5856 5598 5868
rect 6546 5788 6552 5840
rect 6604 5828 6610 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6604 5800 6653 5828
rect 6604 5788 6610 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 6641 5791 6699 5797
rect 2682 5652 2688 5704
rect 2740 5692 2746 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2740 5664 3065 5692
rect 2740 5652 2746 5664
rect 3053 5661 3065 5664
rect 3099 5692 3111 5695
rect 3142 5692 3148 5704
rect 3099 5664 3148 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 6086 5692 6092 5704
rect 5460 5664 6092 5692
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 2869 5627 2927 5633
rect 2869 5624 2881 5627
rect 2648 5596 2881 5624
rect 2648 5584 2654 5596
rect 2869 5593 2881 5596
rect 2915 5593 2927 5627
rect 2869 5587 2927 5593
rect 4985 5627 5043 5633
rect 4985 5593 4997 5627
rect 5031 5593 5043 5627
rect 4985 5587 5043 5593
rect 5169 5627 5227 5633
rect 5169 5593 5181 5627
rect 5215 5624 5227 5627
rect 5460 5624 5488 5664
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6748 5692 6776 5868
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 14090 5856 14096 5908
rect 14148 5856 14154 5908
rect 14921 5899 14979 5905
rect 14921 5865 14933 5899
rect 14967 5896 14979 5899
rect 15286 5896 15292 5908
rect 14967 5868 15292 5896
rect 14967 5865 14979 5868
rect 14921 5859 14979 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 18322 5896 18328 5908
rect 15896 5868 18328 5896
rect 15896 5856 15902 5868
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 21726 5856 21732 5908
rect 21784 5896 21790 5908
rect 22094 5896 22100 5908
rect 21784 5868 22100 5896
rect 21784 5856 21790 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 23106 5856 23112 5908
rect 23164 5896 23170 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 23164 5868 23857 5896
rect 23164 5856 23170 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 23934 5856 23940 5908
rect 23992 5896 23998 5908
rect 25314 5896 25320 5908
rect 23992 5868 25320 5896
rect 23992 5856 23998 5868
rect 25314 5856 25320 5868
rect 25372 5856 25378 5908
rect 25774 5856 25780 5908
rect 25832 5856 25838 5908
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5828 8263 5831
rect 8294 5828 8300 5840
rect 8251 5800 8300 5828
rect 8251 5797 8263 5800
rect 8205 5791 8263 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 13814 5788 13820 5840
rect 13872 5788 13878 5840
rect 14182 5788 14188 5840
rect 14240 5828 14246 5840
rect 14734 5828 14740 5840
rect 14240 5800 14740 5828
rect 14240 5788 14246 5800
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 16942 5788 16948 5840
rect 17000 5828 17006 5840
rect 17218 5828 17224 5840
rect 17000 5800 17224 5828
rect 17000 5788 17006 5800
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 17678 5788 17684 5840
rect 17736 5788 17742 5840
rect 19334 5788 19340 5840
rect 19392 5828 19398 5840
rect 20530 5828 20536 5840
rect 19392 5800 20536 5828
rect 19392 5788 19398 5800
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 23750 5788 23756 5840
rect 23808 5828 23814 5840
rect 25409 5831 25467 5837
rect 25409 5828 25421 5831
rect 23808 5800 25421 5828
rect 23808 5788 23814 5800
rect 25409 5797 25421 5800
rect 25455 5797 25467 5831
rect 25409 5791 25467 5797
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5760 8171 5763
rect 8754 5760 8760 5772
rect 8159 5732 8760 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 7846 5695 7904 5701
rect 7846 5692 7858 5695
rect 6748 5664 7858 5692
rect 7846 5661 7858 5664
rect 7892 5661 7904 5695
rect 8772 5692 8800 5720
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 8772 5664 10333 5692
rect 7846 5655 7904 5661
rect 10321 5661 10333 5664
rect 10367 5692 10379 5695
rect 10502 5692 10508 5704
rect 10367 5664 10508 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10778 5701 10784 5704
rect 10772 5692 10784 5701
rect 10739 5664 10784 5692
rect 10772 5655 10784 5664
rect 10778 5652 10784 5655
rect 10836 5652 10842 5704
rect 13832 5692 13860 5788
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 14056 5732 15332 5760
rect 14056 5720 14062 5732
rect 14384 5701 14412 5732
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13832 5664 13921 5692
rect 13909 5661 13921 5664
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 15102 5652 15108 5704
rect 15160 5652 15166 5704
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 5534 5633 5540 5636
rect 5215 5596 5488 5624
rect 5215 5593 5227 5596
rect 5169 5587 5227 5593
rect 5528 5587 5540 5633
rect 3234 5516 3240 5568
rect 3292 5516 3298 5568
rect 5000 5556 5028 5587
rect 5534 5584 5540 5587
rect 5592 5584 5598 5636
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 7800 5596 8585 5624
rect 7800 5584 7806 5596
rect 8573 5593 8585 5596
rect 8619 5624 8631 5627
rect 9306 5624 9312 5636
rect 8619 5596 9312 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 10054 5627 10112 5633
rect 10054 5624 10066 5627
rect 9548 5596 10066 5624
rect 9548 5584 9554 5596
rect 10054 5593 10066 5596
rect 10100 5593 10112 5627
rect 10054 5587 10112 5593
rect 13725 5627 13783 5633
rect 13725 5593 13737 5627
rect 13771 5624 13783 5627
rect 13814 5624 13820 5636
rect 13771 5596 13820 5624
rect 13771 5593 13783 5596
rect 13725 5587 13783 5593
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 14090 5584 14096 5636
rect 14148 5624 14154 5636
rect 15212 5624 15240 5655
rect 14148 5596 15240 5624
rect 14148 5584 14154 5596
rect 6454 5556 6460 5568
rect 5000 5528 6460 5556
rect 6454 5516 6460 5528
rect 6512 5556 6518 5568
rect 6638 5556 6644 5568
rect 6512 5528 6644 5556
rect 6512 5516 6518 5528
rect 6638 5516 6644 5528
rect 6696 5556 6702 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6696 5528 6745 5556
rect 6696 5516 6702 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8720 5528 8769 5556
rect 8720 5516 8726 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 11974 5556 11980 5568
rect 11931 5528 11980 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 14550 5556 14556 5568
rect 13587 5528 14556 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 15304 5556 15332 5732
rect 15562 5720 15568 5772
rect 15620 5720 15626 5772
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 17770 5760 17776 5772
rect 16816 5732 17776 5760
rect 16816 5720 16822 5732
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 15654 5692 15660 5704
rect 15519 5664 15660 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 17696 5701 17724 5732
rect 17770 5720 17776 5732
rect 17828 5760 17834 5772
rect 17828 5732 18276 5760
rect 17828 5720 17834 5732
rect 18248 5704 18276 5732
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19116 5732 20760 5760
rect 19116 5720 19122 5732
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 17865 5695 17923 5701
rect 17865 5661 17877 5695
rect 17911 5692 17923 5695
rect 17911 5664 18184 5692
rect 17911 5661 17923 5664
rect 17865 5655 17923 5661
rect 15838 5633 15844 5636
rect 15832 5587 15844 5633
rect 15838 5584 15844 5587
rect 15896 5584 15902 5636
rect 17218 5584 17224 5636
rect 17276 5584 17282 5636
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 18049 5627 18107 5633
rect 18049 5624 18061 5627
rect 17460 5596 18061 5624
rect 17460 5584 17466 5596
rect 18049 5593 18061 5596
rect 18095 5593 18107 5627
rect 18156 5624 18184 5664
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18432 5624 18460 5655
rect 20254 5652 20260 5704
rect 20312 5652 20318 5704
rect 20732 5701 20760 5732
rect 24412 5732 25084 5760
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 22186 5692 22192 5704
rect 20763 5664 22192 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 20548 5624 20576 5655
rect 22186 5652 22192 5664
rect 22244 5692 22250 5704
rect 22646 5692 22652 5704
rect 22244 5664 22652 5692
rect 22244 5652 22250 5664
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 23753 5695 23811 5701
rect 23753 5692 23765 5695
rect 23492 5664 23765 5692
rect 18156 5596 20576 5624
rect 18049 5587 18107 5593
rect 16114 5556 16120 5568
rect 15304 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 17034 5516 17040 5568
rect 17092 5516 17098 5568
rect 20548 5556 20576 5596
rect 20625 5627 20683 5633
rect 20625 5593 20637 5627
rect 20671 5624 20683 5627
rect 20806 5624 20812 5636
rect 20671 5596 20812 5624
rect 20671 5593 20683 5596
rect 20625 5587 20683 5593
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 20984 5627 21042 5633
rect 20984 5593 20996 5627
rect 21030 5624 21042 5627
rect 21358 5624 21364 5636
rect 21030 5596 21364 5624
rect 21030 5593 21042 5596
rect 20984 5587 21042 5593
rect 21358 5584 21364 5596
rect 21416 5584 21422 5636
rect 21542 5584 21548 5636
rect 21600 5624 21606 5636
rect 23492 5624 23520 5664
rect 23753 5661 23765 5664
rect 23799 5692 23811 5695
rect 23799 5664 24164 5692
rect 23799 5661 23811 5664
rect 23753 5655 23811 5661
rect 21600 5596 23520 5624
rect 23569 5627 23627 5633
rect 21600 5584 21606 5596
rect 23569 5593 23581 5627
rect 23615 5624 23627 5627
rect 23934 5624 23940 5636
rect 23615 5596 23940 5624
rect 23615 5593 23627 5596
rect 23569 5587 23627 5593
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 24026 5584 24032 5636
rect 24084 5584 24090 5636
rect 24136 5624 24164 5664
rect 24213 5627 24271 5633
rect 24213 5624 24225 5627
rect 24136 5596 24225 5624
rect 24213 5593 24225 5596
rect 24259 5624 24271 5627
rect 24412 5624 24440 5732
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5692 24731 5695
rect 24854 5692 24860 5704
rect 24719 5664 24860 5692
rect 24719 5661 24731 5664
rect 24673 5655 24731 5661
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 25056 5701 25084 5732
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 25041 5695 25099 5701
rect 25041 5661 25053 5695
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 24259 5596 24440 5624
rect 24259 5593 24271 5596
rect 24213 5587 24271 5593
rect 24762 5584 24768 5636
rect 24820 5584 24826 5636
rect 24964 5624 24992 5655
rect 25590 5652 25596 5704
rect 25648 5652 25654 5704
rect 25225 5627 25283 5633
rect 25225 5624 25237 5627
rect 24964 5596 25237 5624
rect 25225 5593 25237 5596
rect 25271 5624 25283 5627
rect 25498 5624 25504 5636
rect 25271 5596 25504 5624
rect 25271 5593 25283 5596
rect 25225 5587 25283 5593
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 21266 5556 21272 5568
rect 20548 5528 21272 5556
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 22094 5516 22100 5568
rect 22152 5556 22158 5568
rect 23290 5556 23296 5568
rect 22152 5528 23296 5556
rect 22152 5516 22158 5528
rect 23290 5516 23296 5528
rect 23348 5516 23354 5568
rect 23385 5559 23443 5565
rect 23385 5525 23397 5559
rect 23431 5556 23443 5559
rect 23474 5556 23480 5568
rect 23431 5528 23480 5556
rect 23431 5525 23443 5528
rect 23385 5519 23443 5525
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 23658 5516 23664 5568
rect 23716 5556 23722 5568
rect 24397 5559 24455 5565
rect 24397 5556 24409 5559
rect 23716 5528 24409 5556
rect 23716 5516 23722 5528
rect 24397 5525 24409 5528
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 1104 5466 26220 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 26220 5466
rect 1104 5392 26220 5414
rect 1946 5312 1952 5364
rect 2004 5312 2010 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 4407 5355 4465 5361
rect 4407 5352 4419 5355
rect 3292 5324 4419 5352
rect 3292 5312 3298 5324
rect 4407 5321 4419 5324
rect 4453 5321 4465 5355
rect 4407 5315 4465 5321
rect 5534 5312 5540 5364
rect 5592 5312 5598 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5810 5352 5816 5364
rect 5767 5324 5816 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 6565 5355 6623 5361
rect 6565 5352 6577 5355
rect 6144 5324 6577 5352
rect 6144 5312 6150 5324
rect 6565 5321 6577 5324
rect 6611 5321 6623 5355
rect 6565 5315 6623 5321
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8570 5352 8576 5364
rect 7883 5324 8576 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 1964 5284 1992 5312
rect 1964 5256 4200 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2682 5216 2688 5228
rect 2179 5188 2688 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 1964 5148 1992 5179
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 4172 5225 4200 5256
rect 4614 5244 4620 5296
rect 4672 5244 4678 5296
rect 6365 5287 6423 5293
rect 6365 5253 6377 5287
rect 6411 5284 6423 5287
rect 6454 5284 6460 5296
rect 6411 5256 6460 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6748 5284 6776 5315
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 14458 5352 14464 5364
rect 13648 5324 14464 5352
rect 7466 5284 7472 5296
rect 6748 5256 7472 5284
rect 3901 5219 3959 5225
rect 3901 5185 3913 5219
rect 3947 5216 3959 5219
rect 4157 5219 4215 5225
rect 3947 5188 4108 5216
rect 3947 5185 3959 5188
rect 3901 5179 3959 5185
rect 4080 5148 4108 5188
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 5258 5216 5264 5228
rect 4203 5188 5264 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5216 6147 5219
rect 6748 5216 6776 5256
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 7653 5287 7711 5293
rect 7653 5253 7665 5287
rect 7699 5284 7711 5287
rect 7926 5284 7932 5296
rect 7699 5256 7932 5284
rect 7699 5253 7711 5256
rect 7653 5247 7711 5253
rect 7926 5244 7932 5256
rect 7984 5244 7990 5296
rect 8754 5244 8760 5296
rect 8812 5284 8818 5296
rect 8812 5256 9352 5284
rect 8812 5244 8818 5256
rect 6135 5188 6776 5216
rect 6135 5185 6147 5188
rect 6089 5179 6147 5185
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 9324 5225 9352 5256
rect 9042 5219 9100 5225
rect 9042 5216 9054 5219
rect 8720 5188 9054 5216
rect 8720 5176 8726 5188
rect 9042 5185 9054 5188
rect 9088 5185 9100 5219
rect 9042 5179 9100 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 13648 5225 13676 5324
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 15838 5352 15844 5364
rect 15795 5324 15844 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19484 5324 19533 5352
rect 19484 5312 19490 5324
rect 19521 5321 19533 5324
rect 19567 5352 19579 5355
rect 19567 5324 20484 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 14001 5287 14059 5293
rect 14001 5284 14013 5287
rect 13740 5256 14013 5284
rect 13740 5225 13768 5256
rect 14001 5253 14013 5256
rect 14047 5253 14059 5287
rect 14001 5247 14059 5253
rect 14369 5287 14427 5293
rect 14369 5253 14381 5287
rect 14415 5284 14427 5287
rect 14642 5284 14648 5296
rect 14415 5256 14648 5284
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 15013 5287 15071 5293
rect 15013 5253 15025 5287
rect 15059 5284 15071 5287
rect 17034 5284 17040 5296
rect 15059 5256 15792 5284
rect 15059 5253 15071 5256
rect 15013 5247 15071 5253
rect 15764 5228 15792 5256
rect 16224 5256 17040 5284
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 13228 5188 13553 5216
rect 13228 5176 13234 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 13556 5148 13584 5179
rect 1964 5120 2636 5148
rect 4080 5120 4292 5148
rect 13556 5120 13676 5148
rect 2608 5092 2636 5120
rect 2041 5083 2099 5089
rect 2041 5049 2053 5083
rect 2087 5080 2099 5083
rect 2409 5083 2467 5089
rect 2087 5052 2360 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 2222 4972 2228 5024
rect 2280 4972 2286 5024
rect 2332 5012 2360 5052
rect 2409 5049 2421 5083
rect 2455 5080 2467 5083
rect 2498 5080 2504 5092
rect 2455 5052 2504 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 4264 5089 4292 5120
rect 2777 5083 2835 5089
rect 2777 5080 2789 5083
rect 2648 5052 2789 5080
rect 2648 5040 2654 5052
rect 2777 5049 2789 5052
rect 2823 5049 2835 5083
rect 2777 5043 2835 5049
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5049 4307 5083
rect 4614 5080 4620 5092
rect 4249 5043 4307 5049
rect 4356 5052 4620 5080
rect 4356 5012 4384 5052
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 7926 5040 7932 5092
rect 7984 5040 7990 5092
rect 2332 4984 4384 5012
rect 4430 4972 4436 5024
rect 4488 4972 4494 5024
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6638 5012 6644 5024
rect 6595 4984 6644 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13648 5012 13676 5120
rect 13924 5080 13952 5179
rect 14090 5176 14096 5228
rect 14148 5216 14154 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 14148 5188 14197 5216
rect 14148 5176 14154 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 15102 5176 15108 5228
rect 15160 5216 15166 5228
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 15160 5188 15209 5216
rect 15160 5176 15166 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15304 5148 15332 5179
rect 15470 5176 15476 5228
rect 15528 5176 15534 5228
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5216 15623 5219
rect 15611 5188 15700 5216
rect 15611 5185 15623 5188
rect 15565 5179 15623 5185
rect 14700 5120 15332 5148
rect 14700 5108 14706 5120
rect 14182 5080 14188 5092
rect 13924 5052 14188 5080
rect 14182 5040 14188 5052
rect 14240 5040 14246 5092
rect 15378 5012 15384 5024
rect 13648 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15672 5012 15700 5188
rect 15746 5176 15752 5228
rect 15804 5176 15810 5228
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16224 5225 16252 5256
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 18230 5244 18236 5296
rect 18288 5284 18294 5296
rect 20349 5287 20407 5293
rect 20349 5284 20361 5287
rect 18288 5256 20361 5284
rect 18288 5244 18294 5256
rect 20349 5253 20361 5256
rect 20395 5253 20407 5287
rect 20349 5247 20407 5253
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 16209 5179 16267 5185
rect 15838 5108 15844 5160
rect 15896 5148 15902 5160
rect 16132 5148 16160 5179
rect 16390 5176 16396 5228
rect 16448 5176 16454 5228
rect 18046 5176 18052 5228
rect 18104 5216 18110 5228
rect 18397 5219 18455 5225
rect 18397 5216 18409 5219
rect 18104 5188 18409 5216
rect 18104 5176 18110 5188
rect 18397 5185 18409 5188
rect 18443 5185 18455 5219
rect 18397 5179 18455 5185
rect 20162 5176 20168 5228
rect 20220 5176 20226 5228
rect 20254 5176 20260 5228
rect 20312 5176 20318 5228
rect 15896 5120 16160 5148
rect 15896 5108 15902 5120
rect 18138 5108 18144 5160
rect 18196 5108 18202 5160
rect 20364 5080 20392 5247
rect 20456 5228 20484 5324
rect 20990 5312 20996 5364
rect 21048 5352 21054 5364
rect 21266 5352 21272 5364
rect 21048 5324 21272 5352
rect 21048 5312 21054 5324
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 22094 5352 22100 5364
rect 21376 5324 22100 5352
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 21376 5284 21404 5324
rect 22094 5312 22100 5324
rect 22152 5312 22158 5364
rect 24029 5355 24087 5361
rect 24029 5321 24041 5355
rect 24075 5352 24087 5355
rect 24075 5324 24256 5352
rect 24075 5321 24087 5324
rect 24029 5315 24087 5321
rect 22186 5284 22192 5296
rect 20864 5256 21404 5284
rect 20864 5244 20870 5256
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20496 5188 20545 5216
rect 20496 5176 20502 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20533 5179 20591 5185
rect 21266 5176 21272 5228
rect 21324 5176 21330 5228
rect 21376 5225 21404 5256
rect 21836 5256 22192 5284
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 21450 5176 21456 5228
rect 21508 5176 21514 5228
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5216 21695 5219
rect 21726 5216 21732 5228
rect 21683 5188 21732 5216
rect 21683 5185 21695 5188
rect 21637 5179 21695 5185
rect 21726 5176 21732 5188
rect 21784 5176 21790 5228
rect 21836 5225 21864 5256
rect 22186 5244 22192 5256
rect 22244 5284 22250 5296
rect 23290 5284 23296 5296
rect 22244 5256 23296 5284
rect 22244 5244 22250 5256
rect 23290 5244 23296 5256
rect 23348 5284 23354 5296
rect 24228 5284 24256 5324
rect 25314 5312 25320 5364
rect 25372 5352 25378 5364
rect 25501 5355 25559 5361
rect 25501 5352 25513 5355
rect 25372 5324 25513 5352
rect 25372 5312 25378 5324
rect 25501 5321 25513 5324
rect 25547 5321 25559 5355
rect 25501 5315 25559 5321
rect 24366 5287 24424 5293
rect 24366 5284 24378 5287
rect 23348 5256 24164 5284
rect 24228 5256 24378 5284
rect 23348 5244 23354 5256
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5185 21879 5219
rect 22077 5219 22135 5225
rect 22077 5216 22089 5219
rect 21821 5179 21879 5185
rect 21928 5188 22089 5216
rect 20993 5151 21051 5157
rect 20993 5117 21005 5151
rect 21039 5148 21051 5151
rect 21928 5148 21956 5188
rect 22077 5185 22089 5188
rect 22123 5185 22135 5219
rect 22077 5179 22135 5185
rect 23014 5176 23020 5228
rect 23072 5216 23078 5228
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 23072 5188 23397 5216
rect 23072 5176 23078 5188
rect 23385 5185 23397 5188
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 23474 5176 23480 5228
rect 23532 5216 23538 5228
rect 23569 5219 23627 5225
rect 23569 5216 23581 5219
rect 23532 5188 23581 5216
rect 23532 5176 23538 5188
rect 23569 5185 23581 5188
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23753 5219 23811 5225
rect 23753 5185 23765 5219
rect 23799 5216 23811 5219
rect 23842 5216 23848 5228
rect 23799 5188 23848 5216
rect 23799 5185 23811 5188
rect 23753 5179 23811 5185
rect 21039 5120 21956 5148
rect 21039 5117 21051 5120
rect 20993 5111 21051 5117
rect 23198 5108 23204 5160
rect 23256 5148 23262 5160
rect 23676 5148 23704 5179
rect 23842 5176 23848 5188
rect 23900 5176 23906 5228
rect 24136 5225 24164 5256
rect 24366 5253 24378 5256
rect 24412 5253 24424 5287
rect 24366 5247 24424 5253
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5185 24179 5219
rect 25516 5216 25544 5315
rect 25774 5312 25780 5364
rect 25832 5312 25838 5364
rect 25593 5219 25651 5225
rect 25593 5216 25605 5219
rect 25516 5188 25605 5216
rect 24121 5179 24179 5185
rect 25593 5185 25605 5188
rect 25639 5185 25651 5219
rect 25593 5179 25651 5185
rect 23256 5120 23888 5148
rect 23256 5108 23262 5120
rect 23860 5092 23888 5120
rect 20530 5080 20536 5092
rect 19904 5052 20116 5080
rect 20364 5052 20536 5080
rect 19904 5012 19932 5052
rect 15672 4984 19932 5012
rect 19978 4972 19984 5024
rect 20036 4972 20042 5024
rect 20088 5012 20116 5052
rect 20530 5040 20536 5052
rect 20588 5040 20594 5092
rect 23658 5080 23664 5092
rect 23124 5052 23664 5080
rect 23124 5012 23152 5052
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 23842 5040 23848 5092
rect 23900 5040 23906 5092
rect 20088 4984 23152 5012
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 1104 4922 26220 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 26220 4922
rect 1104 4848 26220 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3513 4811 3571 4817
rect 3513 4808 3525 4811
rect 2832 4780 3525 4808
rect 2832 4768 2838 4780
rect 3513 4777 3525 4780
rect 3559 4777 3571 4811
rect 3513 4771 3571 4777
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8386 4808 8392 4820
rect 8343 4780 8392 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14642 4808 14648 4820
rect 13872 4780 14648 4808
rect 13872 4768 13878 4780
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 14734 4768 14740 4820
rect 14792 4808 14798 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14792 4780 15117 4808
rect 14792 4768 14798 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15528 4780 15853 4808
rect 15528 4768 15534 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 18874 4768 18880 4820
rect 18932 4768 18938 4820
rect 20990 4808 20996 4820
rect 18984 4780 20996 4808
rect 18322 4740 18328 4752
rect 18248 4712 18328 4740
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 2004 4644 2145 4672
rect 2004 4632 2010 4644
rect 2133 4641 2145 4644
rect 2179 4641 2191 4675
rect 8478 4672 8484 4684
rect 2133 4635 2191 4641
rect 8220 4644 8484 4672
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 8220 4613 8248 4644
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 16758 4672 16764 4684
rect 16040 4644 16764 4672
rect 16040 4616 16068 4644
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 2389 4607 2447 4613
rect 2389 4604 2401 4607
rect 2280 4576 2401 4604
rect 2280 4564 2286 4576
rect 2389 4573 2401 4576
rect 2435 4573 2447 4607
rect 2389 4567 2447 4573
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8352 4576 8401 4604
rect 8352 4564 8358 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 12526 4564 12532 4616
rect 12584 4564 12590 4616
rect 12796 4607 12854 4613
rect 12796 4573 12808 4607
rect 12842 4604 12854 4607
rect 13262 4604 13268 4616
rect 12842 4576 13268 4604
rect 12842 4573 12854 4576
rect 12796 4567 12854 4573
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 14366 4564 14372 4616
rect 14424 4564 14430 4616
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14734 4564 14740 4616
rect 14792 4564 14798 4616
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 14936 4536 14964 4567
rect 16022 4564 16028 4616
rect 16080 4564 16086 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 17954 4604 17960 4616
rect 16439 4576 17960 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18248 4604 18276 4712
rect 18322 4700 18328 4712
rect 18380 4740 18386 4752
rect 18984 4740 19012 4780
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 21450 4768 21456 4820
rect 21508 4808 21514 4820
rect 21637 4811 21695 4817
rect 21637 4808 21649 4811
rect 21508 4780 21649 4808
rect 21508 4768 21514 4780
rect 21637 4777 21649 4780
rect 21683 4777 21695 4811
rect 21637 4771 21695 4777
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21784 4780 21925 4808
rect 21784 4768 21790 4780
rect 21913 4777 21925 4780
rect 21959 4777 21971 4811
rect 21913 4771 21971 4777
rect 25498 4768 25504 4820
rect 25556 4808 25562 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 25556 4780 25789 4808
rect 25556 4768 25562 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 25777 4771 25835 4777
rect 21818 4740 21824 4752
rect 18380 4712 19012 4740
rect 19352 4712 21824 4740
rect 18380 4700 18386 4712
rect 18305 4607 18363 4613
rect 18305 4604 18317 4607
rect 18248 4576 18317 4604
rect 18305 4573 18317 4576
rect 18351 4573 18363 4607
rect 18305 4567 18363 4573
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4573 18567 4607
rect 18509 4567 18567 4573
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 18874 4604 18880 4616
rect 18739 4576 18880 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 12820 4508 14964 4536
rect 12820 4480 12848 4508
rect 12802 4428 12808 4480
rect 12860 4428 12866 4480
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 13998 4468 14004 4480
rect 13955 4440 14004 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14090 4428 14096 4480
rect 14148 4428 14154 4480
rect 14936 4468 14964 4508
rect 16114 4496 16120 4548
rect 16172 4496 16178 4548
rect 16206 4496 16212 4548
rect 16264 4496 16270 4548
rect 17678 4496 17684 4548
rect 17736 4536 17742 4548
rect 18432 4536 18460 4567
rect 17736 4508 18460 4536
rect 18524 4536 18552 4567
rect 18874 4564 18880 4576
rect 18932 4564 18938 4616
rect 18966 4564 18972 4616
rect 19024 4604 19030 4616
rect 19061 4607 19119 4613
rect 19061 4604 19073 4607
rect 19024 4576 19073 4604
rect 19024 4564 19030 4576
rect 19061 4573 19073 4576
rect 19107 4604 19119 4607
rect 19352 4604 19380 4712
rect 21818 4700 21824 4712
rect 21876 4700 21882 4752
rect 23198 4672 23204 4684
rect 21468 4644 23204 4672
rect 19107 4576 19380 4604
rect 19107 4573 19119 4576
rect 19061 4567 19119 4573
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 21468 4613 21496 4644
rect 23198 4632 23204 4644
rect 23256 4632 23262 4684
rect 23290 4632 23296 4684
rect 23348 4672 23354 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23348 4644 24409 4672
rect 23348 4632 23354 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 20312 4576 21465 4604
rect 20312 4564 20318 4576
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 21634 4564 21640 4616
rect 21692 4604 21698 4616
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 21692 4576 21741 4604
rect 21692 4564 21698 4576
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 21729 4567 21787 4573
rect 23014 4564 23020 4616
rect 23072 4604 23078 4616
rect 23569 4607 23627 4613
rect 23569 4604 23581 4607
rect 23072 4576 23581 4604
rect 23072 4564 23078 4576
rect 19245 4539 19303 4545
rect 19245 4536 19257 4539
rect 18524 4508 19257 4536
rect 17736 4496 17742 4508
rect 17034 4468 17040 4480
rect 14936 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 18432 4468 18460 4508
rect 19245 4505 19257 4508
rect 19291 4505 19303 4539
rect 19245 4499 19303 4505
rect 19518 4496 19524 4548
rect 19576 4536 19582 4548
rect 19613 4539 19671 4545
rect 19613 4536 19625 4539
rect 19576 4508 19625 4536
rect 19576 4496 19582 4508
rect 19613 4505 19625 4508
rect 19659 4505 19671 4539
rect 19613 4499 19671 4505
rect 21269 4539 21327 4545
rect 21269 4505 21281 4539
rect 21315 4536 21327 4539
rect 21542 4536 21548 4548
rect 21315 4508 21548 4536
rect 21315 4505 21327 4508
rect 21269 4499 21327 4505
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 19426 4468 19432 4480
rect 18432 4440 19432 4468
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 21726 4428 21732 4480
rect 21784 4468 21790 4480
rect 23032 4468 23060 4564
rect 23308 4548 23336 4576
rect 23569 4573 23581 4576
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 23750 4564 23756 4616
rect 23808 4564 23814 4616
rect 23842 4564 23848 4616
rect 23900 4564 23906 4616
rect 23937 4607 23995 4613
rect 23937 4573 23949 4607
rect 23983 4604 23995 4607
rect 24118 4604 24124 4616
rect 23983 4576 24124 4604
rect 23983 4573 23995 4576
rect 23937 4567 23995 4573
rect 24118 4564 24124 4576
rect 24176 4564 24182 4616
rect 24412 4604 24440 4635
rect 24412 4576 24900 4604
rect 23290 4496 23296 4548
rect 23348 4496 23354 4548
rect 21784 4440 23060 4468
rect 21784 4428 21790 4440
rect 23106 4428 23112 4480
rect 23164 4468 23170 4480
rect 23860 4468 23888 4564
rect 24872 4548 24900 4576
rect 24213 4539 24271 4545
rect 24213 4505 24225 4539
rect 24259 4536 24271 4539
rect 24642 4539 24700 4545
rect 24642 4536 24654 4539
rect 24259 4508 24654 4536
rect 24259 4505 24271 4508
rect 24213 4499 24271 4505
rect 24642 4505 24654 4508
rect 24688 4505 24700 4539
rect 24642 4499 24700 4505
rect 24854 4496 24860 4548
rect 24912 4496 24918 4548
rect 24762 4468 24768 4480
rect 23164 4440 24768 4468
rect 23164 4428 23170 4440
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 1104 4378 26220 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 26220 4378
rect 1104 4304 26220 4326
rect 14734 4224 14740 4276
rect 14792 4224 14798 4276
rect 17402 4264 17408 4276
rect 16684 4236 17408 4264
rect 14752 4196 14780 4224
rect 16684 4205 16712 4236
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 19610 4224 19616 4276
rect 19668 4224 19674 4276
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 21542 4264 21548 4276
rect 20220 4236 20668 4264
rect 20220 4224 20226 4236
rect 16669 4199 16727 4205
rect 14752 4168 16528 4196
rect 12888 4131 12946 4137
rect 12888 4097 12900 4131
rect 12934 4128 12946 4131
rect 14090 4128 14096 4140
rect 12934 4100 14096 4128
rect 12934 4097 12946 4100
rect 12888 4091 12946 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15028 4137 15056 4168
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14424 4100 14657 4128
rect 14424 4088 14430 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4097 14887 4131
rect 14829 4091 14887 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12621 4063 12679 4069
rect 12621 4060 12633 4063
rect 12584 4032 12633 4060
rect 12584 4020 12590 4032
rect 12621 4029 12633 4032
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 12636 3924 12664 4023
rect 14752 3992 14780 4091
rect 14844 4060 14872 4091
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 15286 4060 15292 4072
rect 14844 4032 15292 4060
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 15488 4060 15516 4091
rect 15562 4088 15568 4140
rect 15620 4088 15626 4140
rect 15764 4137 15792 4168
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 15838 4088 15844 4140
rect 15896 4088 15902 4140
rect 16022 4088 16028 4140
rect 16080 4088 16086 4140
rect 16117 4131 16175 4137
rect 16117 4097 16129 4131
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 15856 4060 15884 4088
rect 15488 4032 15884 4060
rect 15488 3992 15516 4032
rect 15930 4020 15936 4072
rect 15988 4060 15994 4072
rect 16132 4060 16160 4091
rect 16206 4088 16212 4140
rect 16264 4088 16270 4140
rect 16390 4088 16396 4140
rect 16448 4088 16454 4140
rect 15988 4032 16160 4060
rect 16500 4060 16528 4168
rect 16669 4165 16681 4199
rect 16715 4165 16727 4199
rect 16669 4159 16727 4165
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 17037 4199 17095 4205
rect 17037 4196 17049 4199
rect 16816 4168 17049 4196
rect 16816 4156 16822 4168
rect 17037 4165 17049 4168
rect 17083 4165 17095 4199
rect 17037 4159 17095 4165
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 19794 4196 19800 4208
rect 18932 4168 19800 4196
rect 18932 4156 18938 4168
rect 19794 4156 19800 4168
rect 19852 4196 19858 4208
rect 19852 4168 20300 4196
rect 19852 4156 19858 4168
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 16942 4128 16948 4140
rect 16899 4100 16948 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4097 17187 4131
rect 17129 4091 17187 4097
rect 17144 4060 17172 4091
rect 17310 4088 17316 4140
rect 17368 4088 17374 4140
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 16500 4032 17172 4060
rect 17420 4060 17448 4091
rect 17494 4088 17500 4140
rect 17552 4088 17558 4140
rect 18138 4088 18144 4140
rect 18196 4088 18202 4140
rect 18408 4131 18466 4137
rect 18408 4097 18420 4131
rect 18454 4128 18466 4131
rect 19242 4128 19248 4140
rect 18454 4100 19248 4128
rect 18454 4097 18466 4100
rect 18408 4091 18466 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 19889 4131 19947 4137
rect 19889 4128 19901 4131
rect 19352 4100 19901 4128
rect 17678 4060 17684 4072
rect 17420 4032 17684 4060
rect 15988 4020 15994 4032
rect 14752 3964 15516 3992
rect 13722 3924 13728 3936
rect 12636 3896 13728 3924
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13872 3896 14013 3924
rect 13872 3884 13878 3896
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 15102 3884 15108 3936
rect 15160 3884 15166 3936
rect 15488 3924 15516 3964
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 15841 3995 15899 4001
rect 15841 3992 15853 3995
rect 15712 3964 15853 3992
rect 15712 3952 15718 3964
rect 15841 3961 15853 3964
rect 15887 3961 15899 3995
rect 16574 3992 16580 4004
rect 15841 3955 15899 3961
rect 16408 3964 16580 3992
rect 16408 3924 16436 3964
rect 16574 3952 16580 3964
rect 16632 3992 16638 4004
rect 17420 3992 17448 4032
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 16632 3964 17448 3992
rect 17696 3964 18184 3992
rect 16632 3952 16638 3964
rect 15488 3896 16436 3924
rect 16482 3884 16488 3936
rect 16540 3924 16546 3936
rect 17696 3924 17724 3964
rect 16540 3896 17724 3924
rect 16540 3884 16546 3896
rect 17770 3884 17776 3936
rect 17828 3884 17834 3936
rect 18156 3924 18184 3964
rect 19352 3924 19380 4100
rect 19889 4097 19901 4100
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 19981 4131 20039 4137
rect 19981 4097 19993 4131
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19996 4060 20024 4091
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 20272 4137 20300 4168
rect 20530 4156 20536 4208
rect 20588 4156 20594 4208
rect 20640 4196 20668 4236
rect 21284 4236 21548 4264
rect 21284 4205 21312 4236
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22554 4264 22560 4276
rect 22152 4236 22560 4264
rect 22152 4224 22158 4236
rect 22554 4224 22560 4236
rect 22612 4264 22618 4276
rect 23014 4264 23020 4276
rect 22612 4236 23020 4264
rect 22612 4224 22618 4236
rect 23014 4224 23020 4236
rect 23072 4224 23078 4276
rect 23106 4224 23112 4276
rect 23164 4224 23170 4276
rect 21269 4199 21327 4205
rect 20640 4168 20760 4196
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20349 4131 20407 4137
rect 20349 4097 20361 4131
rect 20395 4097 20407 4131
rect 20349 4091 20407 4097
rect 19484 4032 20024 4060
rect 19484 4020 19490 4032
rect 19521 3995 19579 4001
rect 19521 3961 19533 3995
rect 19567 3992 19579 3995
rect 19702 3992 19708 4004
rect 19567 3964 19708 3992
rect 19567 3961 19579 3964
rect 19521 3955 19579 3961
rect 19702 3952 19708 3964
rect 19760 3992 19766 4004
rect 20364 3992 20392 4091
rect 20438 4088 20444 4140
rect 20496 4088 20502 4140
rect 20732 4137 20760 4168
rect 21269 4165 21281 4199
rect 21315 4165 21327 4199
rect 21269 4159 21327 4165
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 23124 4196 23152 4224
rect 23566 4196 23572 4208
rect 21508 4168 23152 4196
rect 23216 4168 23572 4196
rect 21508 4156 21514 4168
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4097 20683 4131
rect 20625 4091 20683 4097
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 21358 4128 21364 4140
rect 20763 4100 21364 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 20456 4004 20484 4088
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20640 4060 20668 4091
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 21726 4088 21732 4140
rect 21784 4128 21790 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21784 4100 21833 4128
rect 21784 4088 21790 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21821 4091 21879 4097
rect 21928 4100 22017 4128
rect 21637 4063 21695 4069
rect 20588 4032 20668 4060
rect 20824 4032 21496 4060
rect 20588 4020 20594 4032
rect 19760 3964 20392 3992
rect 19760 3952 19766 3964
rect 20438 3952 20444 4004
rect 20496 3952 20502 4004
rect 20824 3924 20852 4032
rect 21468 3992 21496 4032
rect 21637 4029 21649 4063
rect 21683 4060 21695 4063
rect 21928 4060 21956 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22094 4088 22100 4140
rect 22152 4088 22158 4140
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 21683 4032 21956 4060
rect 21683 4029 21695 4032
rect 21637 4023 21695 4029
rect 22204 3992 22232 4091
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22888 4100 22937 4128
rect 22888 4088 22894 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 23014 4088 23020 4140
rect 23072 4088 23078 4140
rect 23109 4131 23167 4137
rect 23109 4097 23121 4131
rect 23155 4128 23167 4131
rect 23216 4128 23244 4168
rect 23566 4156 23572 4168
rect 23624 4156 23630 4208
rect 24504 4168 24992 4196
rect 23155 4100 23244 4128
rect 23155 4097 23167 4100
rect 23109 4091 23167 4097
rect 23290 4088 23296 4140
rect 23348 4088 23354 4140
rect 24504 4128 24532 4168
rect 23400 4100 24532 4128
rect 24601 4131 24659 4137
rect 22278 4020 22284 4072
rect 22336 4060 22342 4072
rect 23400 4060 23428 4100
rect 24601 4097 24613 4131
rect 24647 4128 24659 4131
rect 24762 4128 24768 4140
rect 24647 4100 24768 4128
rect 24647 4097 24659 4100
rect 24601 4091 24659 4097
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 24854 4088 24860 4140
rect 24912 4088 24918 4140
rect 24964 4128 24992 4168
rect 25225 4131 25283 4137
rect 25225 4128 25237 4131
rect 24964 4100 25237 4128
rect 25225 4097 25237 4100
rect 25271 4097 25283 4131
rect 25225 4091 25283 4097
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 25593 4131 25651 4137
rect 25593 4128 25605 4131
rect 25556 4100 25605 4128
rect 25556 4088 25562 4100
rect 25593 4097 25605 4100
rect 25639 4097 25651 4131
rect 25593 4091 25651 4097
rect 22336 4032 23428 4060
rect 22336 4020 22342 4032
rect 21468 3964 22232 3992
rect 25406 3952 25412 4004
rect 25464 3952 25470 4004
rect 25774 3952 25780 4004
rect 25832 3952 25838 4004
rect 18156 3896 20852 3924
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3924 20959 3927
rect 21174 3924 21180 3936
rect 20947 3896 21180 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 22462 3884 22468 3936
rect 22520 3884 22526 3936
rect 22649 3927 22707 3933
rect 22649 3893 22661 3927
rect 22695 3924 22707 3927
rect 22922 3924 22928 3936
rect 22695 3896 22928 3924
rect 22695 3893 22707 3896
rect 22649 3887 22707 3893
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23106 3884 23112 3936
rect 23164 3924 23170 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 23164 3896 23489 3924
rect 23164 3884 23170 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 23477 3887 23535 3893
rect 1104 3834 26220 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 26220 3834
rect 1104 3760 26220 3782
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 16114 3720 16120 3732
rect 15519 3692 16120 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16540 3692 18644 3720
rect 16540 3680 16546 3692
rect 18616 3584 18644 3692
rect 18966 3680 18972 3732
rect 19024 3680 19030 3732
rect 19242 3680 19248 3732
rect 19300 3680 19306 3732
rect 23106 3720 23112 3732
rect 20180 3692 23112 3720
rect 18690 3612 18696 3664
rect 18748 3652 18754 3664
rect 18748 3624 19932 3652
rect 18748 3612 18754 3624
rect 19334 3584 19340 3596
rect 18616 3556 19340 3584
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 19484 3556 19656 3584
rect 19484 3544 19490 3556
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13780 3488 14105 3516
rect 13780 3476 13786 3488
rect 14093 3485 14105 3488
rect 14139 3516 14151 3519
rect 15470 3516 15476 3528
rect 14139 3488 15476 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 15470 3476 15476 3488
rect 15528 3516 15534 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15528 3488 15853 3516
rect 15528 3476 15534 3488
rect 15841 3485 15853 3488
rect 15887 3516 15899 3519
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 15887 3488 17325 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 17313 3485 17325 3488
rect 17359 3516 17371 3519
rect 18138 3516 18144 3528
rect 17359 3488 18144 3516
rect 17359 3485 17371 3488
rect 17313 3479 17371 3485
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 19628 3525 19656 3556
rect 19794 3544 19800 3596
rect 19852 3544 19858 3596
rect 19904 3584 19932 3624
rect 20180 3584 20208 3692
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 23566 3680 23572 3732
rect 23624 3720 23630 3732
rect 23661 3723 23719 3729
rect 23661 3720 23673 3723
rect 23624 3692 23673 3720
rect 23624 3680 23630 3692
rect 23661 3689 23673 3692
rect 23707 3689 23719 3723
rect 23661 3683 23719 3689
rect 24762 3680 24768 3732
rect 24820 3720 24826 3732
rect 25041 3723 25099 3729
rect 25041 3720 25053 3723
rect 24820 3692 25053 3720
rect 24820 3680 24826 3692
rect 25041 3689 25053 3692
rect 25087 3689 25099 3723
rect 25041 3683 25099 3689
rect 23382 3612 23388 3664
rect 23440 3652 23446 3664
rect 23440 3624 25636 3652
rect 23440 3612 23446 3624
rect 22097 3587 22155 3593
rect 19904 3556 20024 3584
rect 20180 3556 20300 3584
rect 19521 3519 19579 3525
rect 19521 3516 19533 3519
rect 19352 3488 19533 3516
rect 19352 3460 19380 3488
rect 19521 3485 19533 3488
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 19702 3476 19708 3528
rect 19760 3476 19766 3528
rect 19812 3513 19840 3544
rect 19996 3525 20024 3556
rect 19889 3519 19947 3525
rect 19889 3513 19901 3519
rect 19812 3485 19901 3513
rect 19935 3485 19947 3519
rect 19889 3479 19947 3485
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 20162 3476 20168 3528
rect 20220 3476 20226 3528
rect 20272 3525 20300 3556
rect 22097 3553 22109 3587
rect 22143 3584 22155 3587
rect 22186 3584 22192 3596
rect 22143 3556 22192 3584
rect 22143 3553 22155 3556
rect 22097 3547 22155 3553
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 23532 3556 24808 3584
rect 23532 3544 23538 3556
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20373 3519 20431 3525
rect 20373 3516 20385 3519
rect 20257 3479 20315 3485
rect 20364 3485 20385 3516
rect 20419 3485 20431 3519
rect 20364 3479 20431 3485
rect 14366 3457 14372 3460
rect 14360 3448 14372 3457
rect 14327 3420 14372 3448
rect 14360 3411 14372 3420
rect 14366 3408 14372 3411
rect 14424 3408 14430 3460
rect 16108 3451 16166 3457
rect 16108 3417 16120 3451
rect 16154 3448 16166 3451
rect 16666 3448 16672 3460
rect 16154 3420 16672 3448
rect 16154 3417 16166 3420
rect 16108 3411 16166 3417
rect 16666 3408 16672 3420
rect 16724 3408 16730 3460
rect 17580 3451 17638 3457
rect 17580 3417 17592 3451
rect 17626 3448 17638 3451
rect 17770 3448 17776 3460
rect 17626 3420 17776 3448
rect 17626 3417 17638 3420
rect 17580 3411 17638 3417
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 18782 3408 18788 3460
rect 18840 3448 18846 3460
rect 18877 3451 18935 3457
rect 18877 3448 18889 3451
rect 18840 3420 18889 3448
rect 18840 3408 18846 3420
rect 18877 3417 18889 3420
rect 18923 3417 18935 3451
rect 18877 3411 18935 3417
rect 19334 3408 19340 3460
rect 19392 3408 19398 3460
rect 20364 3448 20392 3479
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20588 3488 21312 3516
rect 20588 3476 20594 3488
rect 20272 3420 20392 3448
rect 20272 3392 20300 3420
rect 16942 3340 16948 3392
rect 17000 3380 17006 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 17000 3352 17233 3380
rect 17000 3340 17006 3352
rect 17221 3349 17233 3352
rect 17267 3380 17279 3383
rect 17678 3380 17684 3392
rect 17267 3352 17684 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 17678 3340 17684 3352
rect 17736 3380 17742 3392
rect 19426 3380 19432 3392
rect 17736 3352 19432 3380
rect 17736 3340 17742 3352
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 20254 3340 20260 3392
rect 20312 3340 20318 3392
rect 20346 3340 20352 3392
rect 20404 3380 20410 3392
rect 20533 3383 20591 3389
rect 20533 3380 20545 3383
rect 20404 3352 20545 3380
rect 20404 3340 20410 3352
rect 20533 3349 20545 3352
rect 20579 3349 20591 3383
rect 20533 3343 20591 3349
rect 20717 3383 20775 3389
rect 20717 3349 20729 3383
rect 20763 3380 20775 3383
rect 21174 3380 21180 3392
rect 20763 3352 21180 3380
rect 20763 3349 20775 3352
rect 20717 3343 20775 3349
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 21284 3380 21312 3488
rect 21542 3476 21548 3528
rect 21600 3516 21606 3528
rect 22462 3525 22468 3528
rect 22456 3516 22468 3525
rect 21600 3488 22094 3516
rect 22423 3488 22468 3516
rect 21600 3476 21606 3488
rect 21818 3408 21824 3460
rect 21876 3457 21882 3460
rect 21876 3411 21888 3457
rect 22066 3448 22094 3488
rect 22456 3479 22468 3488
rect 22462 3476 22468 3479
rect 22520 3476 22526 3528
rect 24029 3519 24087 3525
rect 24029 3516 24041 3519
rect 23400 3488 24041 3516
rect 23400 3448 23428 3488
rect 24029 3485 24041 3488
rect 24075 3516 24087 3519
rect 24118 3516 24124 3528
rect 24075 3488 24124 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 24397 3519 24455 3525
rect 24397 3485 24409 3519
rect 24443 3485 24455 3519
rect 24397 3479 24455 3485
rect 22066 3420 23428 3448
rect 21876 3408 21882 3411
rect 23474 3408 23480 3460
rect 23532 3448 23538 3460
rect 23532 3420 23796 3448
rect 23532 3408 23538 3420
rect 22830 3380 22836 3392
rect 21284 3352 22836 3380
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 23569 3383 23627 3389
rect 23569 3380 23581 3383
rect 23072 3352 23581 3380
rect 23072 3340 23078 3352
rect 23569 3349 23581 3352
rect 23615 3349 23627 3383
rect 23768 3380 23796 3420
rect 23842 3408 23848 3460
rect 23900 3408 23906 3460
rect 24412 3380 24440 3479
rect 24486 3476 24492 3528
rect 24544 3516 24550 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24544 3488 24593 3516
rect 24544 3476 24550 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24670 3476 24676 3528
rect 24728 3476 24734 3528
rect 24780 3525 24808 3556
rect 25608 3525 25636 3624
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 25593 3519 25651 3525
rect 25593 3485 25605 3519
rect 25639 3485 25651 3519
rect 25593 3479 25651 3485
rect 23768 3352 24440 3380
rect 23569 3343 23627 3349
rect 25774 3340 25780 3392
rect 25832 3340 25838 3392
rect 1104 3290 26220 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 26220 3290
rect 1104 3216 26220 3238
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15562 3176 15568 3188
rect 15243 3148 15568 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 16666 3136 16672 3188
rect 16724 3136 16730 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 16816 3148 17172 3176
rect 16816 3136 16822 3148
rect 13992 3111 14050 3117
rect 13992 3077 14004 3111
rect 14038 3108 14050 3111
rect 15102 3108 15108 3120
rect 14038 3080 15108 3108
rect 14038 3077 14050 3080
rect 13992 3071 14050 3077
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15657 3111 15715 3117
rect 15657 3108 15669 3111
rect 15344 3080 15669 3108
rect 15344 3068 15350 3080
rect 15657 3077 15669 3080
rect 15703 3077 15715 3111
rect 15657 3071 15715 3077
rect 15841 3111 15899 3117
rect 15841 3077 15853 3111
rect 15887 3108 15899 3111
rect 16114 3108 16120 3120
rect 15887 3080 16120 3108
rect 15887 3077 15899 3080
rect 15841 3071 15899 3077
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 16632 3080 17080 3108
rect 16632 3068 16638 3080
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 15392 3043 15450 3049
rect 15392 3009 15404 3043
rect 15438 3040 15450 3043
rect 15565 3043 15623 3049
rect 15438 3012 15507 3040
rect 15438 3009 15450 3012
rect 15392 3003 15450 3009
rect 15479 2972 15507 3012
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15611 3012 16037 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 15930 2972 15936 2984
rect 15479 2944 15936 2972
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 15194 2904 15200 2916
rect 15151 2876 15200 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 15194 2864 15200 2876
rect 15252 2904 15258 2916
rect 15479 2904 15507 2944
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16040 2972 16068 3003
rect 16942 3000 16948 3052
rect 17000 3000 17006 3052
rect 17052 3049 17080 3080
rect 17144 3049 17172 3148
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 17368 3148 17509 3176
rect 17368 3136 17374 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 19610 3176 19616 3188
rect 17497 3139 17555 3145
rect 19260 3148 19616 3176
rect 17681 3111 17739 3117
rect 17681 3077 17693 3111
rect 17727 3108 17739 3111
rect 18322 3108 18328 3120
rect 17727 3080 18328 3108
rect 17727 3077 17739 3080
rect 17681 3071 17739 3077
rect 18322 3068 18328 3080
rect 18380 3108 18386 3120
rect 18690 3108 18696 3120
rect 18380 3080 18696 3108
rect 18380 3068 18386 3080
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 19092 3111 19150 3117
rect 19092 3077 19104 3111
rect 19138 3108 19150 3111
rect 19260 3108 19288 3148
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 19794 3136 19800 3188
rect 19852 3136 19858 3188
rect 19886 3136 19892 3188
rect 19944 3176 19950 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 19944 3148 20269 3176
rect 19944 3136 19950 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 20346 3136 20352 3188
rect 20404 3176 20410 3188
rect 20404 3148 20852 3176
rect 20404 3136 20410 3148
rect 19138 3080 19288 3108
rect 20272 3080 20484 3108
rect 19138 3077 19150 3080
rect 19092 3071 19150 3077
rect 20272 3052 20300 3080
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 17310 3000 17316 3052
rect 17368 3000 17374 3052
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 17862 3040 17868 3052
rect 17460 3012 17868 3040
rect 17460 3000 17466 3012
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 18782 3040 18788 3052
rect 18340 3012 18788 3040
rect 17420 2972 17448 3000
rect 16040 2944 17448 2972
rect 15252 2876 15507 2904
rect 15252 2864 15258 2876
rect 17034 2864 17040 2916
rect 17092 2904 17098 2916
rect 17310 2904 17316 2916
rect 17092 2876 17316 2904
rect 17092 2864 17098 2876
rect 17310 2864 17316 2876
rect 17368 2904 17374 2916
rect 18340 2904 18368 3012
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 19518 3040 19524 3052
rect 19475 3012 19524 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 19702 3040 19708 3052
rect 19659 3012 19708 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 20254 3000 20260 3052
rect 20312 3000 20318 3052
rect 20456 3049 20484 3080
rect 20622 3068 20628 3120
rect 20680 3068 20686 3120
rect 20824 3049 20852 3148
rect 21082 3136 21088 3188
rect 21140 3176 21146 3188
rect 21453 3179 21511 3185
rect 21453 3176 21465 3179
rect 21140 3148 21465 3176
rect 21140 3136 21146 3148
rect 21453 3145 21465 3148
rect 21499 3145 21511 3179
rect 21453 3139 21511 3145
rect 21818 3136 21824 3188
rect 21876 3136 21882 3188
rect 22186 3176 22192 3188
rect 22066 3148 22192 3176
rect 20990 3068 20996 3120
rect 21048 3108 21054 3120
rect 22066 3108 22094 3148
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 22462 3136 22468 3188
rect 22520 3176 22526 3188
rect 23290 3176 23296 3188
rect 22520 3148 23296 3176
rect 22520 3136 22526 3148
rect 23290 3136 23296 3148
rect 23348 3136 23354 3188
rect 23842 3136 23848 3188
rect 23900 3176 23906 3188
rect 24029 3179 24087 3185
rect 24029 3176 24041 3179
rect 23900 3148 24041 3176
rect 23900 3136 23906 3148
rect 24029 3145 24041 3148
rect 24075 3145 24087 3179
rect 24029 3139 24087 3145
rect 24486 3136 24492 3188
rect 24544 3136 24550 3188
rect 22922 3117 22928 3120
rect 22916 3108 22928 3117
rect 21048 3080 22692 3108
rect 22883 3080 22928 3108
rect 21048 3068 21054 3080
rect 20417 3043 20484 3049
rect 20417 3009 20429 3043
rect 20463 3012 20484 3043
rect 20533 3043 20591 3049
rect 20463 3009 20475 3012
rect 20417 3003 20475 3009
rect 20533 3009 20545 3043
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 17368 2876 18368 2904
rect 19352 2904 19380 2935
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 20548 2972 20576 3003
rect 20898 3000 20904 3052
rect 20956 3000 20962 3052
rect 21082 3000 21088 3052
rect 21140 3000 21146 3052
rect 21174 3000 21180 3052
rect 21232 3000 21238 3052
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21358 3040 21364 3052
rect 21315 3012 21364 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 22094 3000 22100 3052
rect 22152 3000 22158 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 20220 2944 20576 2972
rect 22204 2972 22232 3003
rect 22278 3000 22284 3052
rect 22336 3000 22342 3052
rect 22462 3000 22468 3052
rect 22520 3000 22526 3052
rect 22664 3049 22692 3080
rect 22916 3071 22928 3080
rect 22922 3068 22928 3071
rect 22980 3068 22986 3120
rect 23106 3068 23112 3120
rect 23164 3068 23170 3120
rect 24118 3068 24124 3120
rect 24176 3068 24182 3120
rect 22649 3043 22707 3049
rect 22649 3009 22661 3043
rect 22695 3009 22707 3043
rect 23124 3040 23152 3068
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 23124 3012 24317 3040
rect 22649 3003 22707 3009
rect 24305 3009 24317 3012
rect 24351 3040 24363 3043
rect 24854 3040 24860 3052
rect 24351 3012 24860 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 24854 3000 24860 3012
rect 24912 3000 24918 3052
rect 25222 3000 25228 3052
rect 25280 3040 25286 3052
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 25280 3012 25605 3040
rect 25280 3000 25286 3012
rect 25593 3009 25605 3012
rect 25639 3009 25651 3043
rect 25593 3003 25651 3009
rect 22554 2972 22560 2984
rect 22204 2944 22560 2972
rect 20220 2932 20226 2944
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 19352 2876 20760 2904
rect 17368 2864 17374 2876
rect 17957 2839 18015 2845
rect 17957 2805 17969 2839
rect 18003 2836 18015 2839
rect 18598 2836 18604 2848
rect 18003 2808 18604 2836
rect 18003 2805 18015 2808
rect 17957 2799 18015 2805
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 19886 2836 19892 2848
rect 19392 2808 19892 2836
rect 19392 2796 19398 2808
rect 19886 2796 19892 2808
rect 19944 2836 19950 2848
rect 20530 2836 20536 2848
rect 19944 2808 20536 2836
rect 19944 2796 19950 2808
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 20732 2836 20760 2876
rect 20990 2836 20996 2848
rect 20732 2808 20996 2836
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21542 2836 21548 2848
rect 21140 2808 21548 2836
rect 21140 2796 21146 2808
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 25774 2796 25780 2848
rect 25832 2796 25838 2848
rect 1104 2746 26220 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 26220 2746
rect 1104 2672 26220 2694
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10468 2604 10609 2632
rect 10468 2592 10474 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 18656 2604 19564 2632
rect 18656 2592 18662 2604
rect 18690 2524 18696 2576
rect 18748 2564 18754 2576
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 18748 2536 19349 2564
rect 18748 2524 18754 2536
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19337 2527 19395 2533
rect 12618 2456 12624 2508
rect 12676 2456 12682 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 19426 2496 19432 2508
rect 18012 2468 19432 2496
rect 18012 2456 18018 2468
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10376 2400 10425 2428
rect 10376 2388 10382 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12308 2400 12357 2428
rect 12308 2388 12314 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 13814 2428 13820 2440
rect 13587 2400 13820 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 13906 2388 13912 2440
rect 13964 2388 13970 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14056 2400 14565 2428
rect 14056 2388 14062 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 16114 2428 16120 2440
rect 15887 2400 16120 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 16850 2428 16856 2440
rect 16531 2400 16856 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17218 2428 17224 2440
rect 17175 2400 17224 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 18322 2388 18328 2440
rect 18380 2388 18386 2440
rect 18432 2437 18460 2468
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 19536 2496 19564 2604
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21324 2604 22017 2632
rect 21324 2592 21330 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 20346 2524 20352 2576
rect 20404 2524 20410 2576
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 22278 2564 22284 2576
rect 21591 2536 22284 2564
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 22278 2524 22284 2536
rect 22336 2524 22342 2576
rect 22373 2567 22431 2573
rect 22373 2533 22385 2567
rect 22419 2533 22431 2567
rect 22373 2527 22431 2533
rect 20364 2496 20392 2524
rect 19536 2468 20392 2496
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 18463 2400 18497 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 18598 2388 18604 2440
rect 18656 2388 18662 2440
rect 19536 2437 19564 2468
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 22388 2496 22416 2527
rect 20956 2468 21864 2496
rect 20956 2456 20962 2468
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 19889 2431 19947 2437
rect 19889 2428 19901 2431
rect 19760 2400 19901 2428
rect 19760 2388 19766 2400
rect 19889 2397 19901 2400
rect 19935 2397 19947 2431
rect 19889 2391 19947 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20438 2428 20444 2440
rect 20395 2400 20444 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 21836 2437 21864 2468
rect 22066 2468 22416 2496
rect 21177 2431 21235 2437
rect 21177 2428 21189 2431
rect 21140 2400 21189 2428
rect 21140 2388 21146 2400
rect 21177 2397 21189 2400
rect 21223 2397 21235 2431
rect 21177 2391 21235 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22066 2428 22094 2468
rect 21968 2400 22094 2428
rect 22189 2431 22247 2437
rect 21968 2388 21974 2400
rect 22189 2397 22201 2431
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23014 2428 23020 2440
rect 22971 2400 23020 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 18785 2363 18843 2369
rect 18785 2329 18797 2363
rect 18831 2360 18843 2363
rect 20070 2360 20076 2372
rect 18831 2332 20076 2360
rect 18831 2329 18843 2332
rect 18785 2323 18843 2329
rect 20070 2320 20076 2332
rect 20128 2320 20134 2372
rect 21361 2363 21419 2369
rect 21361 2360 21373 2363
rect 21192 2332 21373 2360
rect 21192 2304 21220 2332
rect 21361 2329 21373 2332
rect 21407 2360 21419 2363
rect 22204 2360 22232 2391
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23256 2400 23305 2428
rect 23256 2388 23262 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23900 2400 23949 2428
rect 23900 2388 23906 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 24854 2388 24860 2440
rect 24912 2388 24918 2440
rect 21407 2332 22232 2360
rect 21407 2329 21419 2332
rect 21361 2323 21419 2329
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 12952 2264 13369 2292
rect 12952 2252 12958 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13596 2264 13737 2292
rect 13596 2252 13602 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 14240 2264 14381 2292
rect 14240 2252 14246 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 14826 2252 14832 2304
rect 14884 2292 14890 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14884 2264 15025 2292
rect 14884 2252 14890 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15528 2264 15669 2292
rect 15528 2252 15534 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16172 2264 16313 2292
rect 16172 2252 16178 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16816 2264 16957 2292
rect 16816 2252 16822 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17460 2264 17601 2292
rect 17460 2252 17466 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 18104 2264 18153 2292
rect 18104 2252 18110 2264
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 19426 2252 19432 2304
rect 19484 2292 19490 2304
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 19484 2264 19717 2292
rect 19484 2252 19490 2264
rect 19705 2261 19717 2264
rect 19751 2261 19763 2295
rect 19705 2255 19763 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20036 2264 20177 2292
rect 20036 2252 20042 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 21174 2252 21180 2304
rect 21232 2252 21238 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22741 2295 22799 2301
rect 22741 2292 22753 2295
rect 22612 2264 22753 2292
rect 22612 2252 22618 2264
rect 22741 2261 22753 2264
rect 22787 2261 22799 2295
rect 22741 2255 22799 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24121 2295 24179 2301
rect 24121 2292 24133 2295
rect 23900 2264 24133 2292
rect 23900 2252 23906 2264
rect 24121 2261 24133 2264
rect 24167 2261 24179 2295
rect 24121 2255 24179 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 24673 2295 24731 2301
rect 24673 2292 24685 2295
rect 24544 2264 24685 2292
rect 24544 2252 24550 2264
rect 24673 2261 24685 2264
rect 24719 2261 24731 2295
rect 24673 2255 24731 2261
rect 1104 2202 26220 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 26220 2202
rect 1104 2128 26220 2150
<< via1 >>
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 12900 27072 12952 27124
rect 13176 26936 13228 26988
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 9404 24760 9456 24812
rect 11888 24760 11940 24812
rect 12072 24803 12124 24812
rect 12072 24769 12106 24803
rect 12106 24769 12124 24803
rect 12072 24760 12124 24769
rect 13912 24760 13964 24812
rect 21732 24760 21784 24812
rect 11796 24735 11848 24744
rect 11796 24701 11805 24735
rect 11805 24701 11839 24735
rect 11839 24701 11848 24735
rect 11796 24692 11848 24701
rect 13360 24692 13412 24744
rect 10876 24624 10928 24676
rect 13176 24667 13228 24676
rect 13176 24633 13185 24667
rect 13185 24633 13219 24667
rect 13219 24633 13228 24667
rect 13176 24624 13228 24633
rect 11060 24599 11112 24608
rect 11060 24565 11069 24599
rect 11069 24565 11103 24599
rect 11103 24565 11112 24599
rect 11060 24556 11112 24565
rect 13268 24599 13320 24608
rect 13268 24565 13277 24599
rect 13277 24565 13311 24599
rect 13311 24565 13320 24599
rect 13268 24556 13320 24565
rect 14280 24599 14332 24608
rect 14280 24565 14289 24599
rect 14289 24565 14323 24599
rect 14323 24565 14332 24599
rect 14280 24556 14332 24565
rect 21180 24599 21232 24608
rect 21180 24565 21189 24599
rect 21189 24565 21223 24599
rect 21223 24565 21232 24599
rect 21180 24556 21232 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 11428 24148 11480 24200
rect 11704 24148 11756 24200
rect 13268 24352 13320 24404
rect 12532 24284 12584 24336
rect 11888 24080 11940 24132
rect 12348 24148 12400 24200
rect 10968 24012 11020 24064
rect 12256 24012 12308 24064
rect 13176 24080 13228 24132
rect 17592 24148 17644 24200
rect 18144 24191 18196 24200
rect 18144 24157 18153 24191
rect 18153 24157 18187 24191
rect 18187 24157 18196 24191
rect 18144 24148 18196 24157
rect 18328 24080 18380 24132
rect 13360 24012 13412 24064
rect 14464 24055 14516 24064
rect 14464 24021 14473 24055
rect 14473 24021 14507 24055
rect 14507 24021 14516 24055
rect 14464 24012 14516 24021
rect 16580 24012 16632 24064
rect 16764 24055 16816 24064
rect 16764 24021 16773 24055
rect 16773 24021 16807 24055
rect 16807 24021 16816 24055
rect 16764 24012 16816 24021
rect 17868 24012 17920 24064
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 19248 24216 19300 24268
rect 19708 24148 19760 24200
rect 23388 24148 23440 24200
rect 19616 24080 19668 24132
rect 21088 24080 21140 24132
rect 21456 24080 21508 24132
rect 19432 24012 19484 24064
rect 20168 24055 20220 24064
rect 20168 24021 20177 24055
rect 20177 24021 20211 24055
rect 20211 24021 20220 24055
rect 20168 24012 20220 24021
rect 21732 24012 21784 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 9404 23851 9456 23860
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 11796 23808 11848 23860
rect 11888 23808 11940 23860
rect 12440 23808 12492 23860
rect 21456 23808 21508 23860
rect 10508 23715 10560 23724
rect 10508 23681 10526 23715
rect 10526 23681 10560 23715
rect 10508 23672 10560 23681
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 10968 23715 11020 23724
rect 10968 23681 10977 23715
rect 10977 23681 11011 23715
rect 11011 23681 11020 23715
rect 10968 23672 11020 23681
rect 12348 23740 12400 23792
rect 14464 23740 14516 23792
rect 16488 23740 16540 23792
rect 12164 23672 12216 23724
rect 12532 23672 12584 23724
rect 14004 23672 14056 23724
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 14740 23715 14792 23724
rect 14740 23681 14749 23715
rect 14749 23681 14783 23715
rect 14783 23681 14792 23715
rect 14740 23672 14792 23681
rect 17960 23672 18012 23724
rect 18144 23740 18196 23792
rect 19156 23672 19208 23724
rect 20628 23672 20680 23724
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 4620 23536 4672 23588
rect 5172 23647 5224 23656
rect 5172 23613 5181 23647
rect 5181 23613 5215 23647
rect 5215 23613 5224 23647
rect 5172 23604 5224 23613
rect 5264 23647 5316 23656
rect 5264 23613 5273 23647
rect 5273 23613 5307 23647
rect 5307 23613 5316 23647
rect 5264 23604 5316 23613
rect 6000 23604 6052 23656
rect 11152 23647 11204 23656
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 11244 23647 11296 23656
rect 11244 23613 11253 23647
rect 11253 23613 11287 23647
rect 11287 23613 11296 23647
rect 11244 23604 11296 23613
rect 13360 23604 13412 23656
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 16212 23647 16264 23656
rect 16212 23613 16221 23647
rect 16221 23613 16255 23647
rect 16255 23613 16264 23647
rect 16212 23604 16264 23613
rect 5448 23468 5500 23520
rect 5540 23511 5592 23520
rect 5540 23477 5549 23511
rect 5549 23477 5583 23511
rect 5583 23477 5592 23511
rect 5540 23468 5592 23477
rect 8668 23511 8720 23520
rect 8668 23477 8677 23511
rect 8677 23477 8711 23511
rect 8711 23477 8720 23511
rect 8668 23468 8720 23477
rect 11336 23511 11388 23520
rect 11336 23477 11345 23511
rect 11345 23477 11379 23511
rect 11379 23477 11388 23511
rect 11336 23468 11388 23477
rect 12992 23511 13044 23520
rect 12992 23477 13001 23511
rect 13001 23477 13035 23511
rect 13035 23477 13044 23511
rect 12992 23468 13044 23477
rect 13084 23468 13136 23520
rect 13820 23468 13872 23520
rect 15568 23468 15620 23520
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 17776 23468 17828 23520
rect 21180 23604 21232 23656
rect 18696 23468 18748 23520
rect 20260 23468 20312 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 3608 23239 3660 23248
rect 3608 23205 3617 23239
rect 3617 23205 3651 23239
rect 3651 23205 3660 23239
rect 3608 23196 3660 23205
rect 3700 23196 3752 23248
rect 5264 23264 5316 23316
rect 8484 23264 8536 23316
rect 10508 23307 10560 23316
rect 10508 23273 10517 23307
rect 10517 23273 10551 23307
rect 10551 23273 10560 23307
rect 10508 23264 10560 23273
rect 3240 23128 3292 23180
rect 4436 23128 4488 23180
rect 4712 23171 4764 23180
rect 4712 23137 4746 23171
rect 4746 23137 4764 23171
rect 4712 23128 4764 23137
rect 10876 23128 10928 23180
rect 1952 23060 2004 23112
rect 5540 23060 5592 23112
rect 8300 23060 8352 23112
rect 11704 23264 11756 23316
rect 11980 23264 12032 23316
rect 12164 23307 12216 23316
rect 12164 23273 12173 23307
rect 12173 23273 12207 23307
rect 12207 23273 12216 23307
rect 12164 23264 12216 23273
rect 12440 23264 12492 23316
rect 13728 23264 13780 23316
rect 14004 23264 14056 23316
rect 16764 23264 16816 23316
rect 11428 23196 11480 23248
rect 11612 23196 11664 23248
rect 12072 23196 12124 23248
rect 14648 23196 14700 23248
rect 11336 23128 11388 23180
rect 2504 23035 2556 23044
rect 2504 23001 2538 23035
rect 2538 23001 2556 23035
rect 2504 22992 2556 23001
rect 4620 22992 4672 23044
rect 2596 22924 2648 22976
rect 5172 22992 5224 23044
rect 7012 22992 7064 23044
rect 8760 22992 8812 23044
rect 11060 23035 11112 23044
rect 11060 23001 11069 23035
rect 11069 23001 11103 23035
rect 11103 23001 11112 23035
rect 11060 22992 11112 23001
rect 11152 23035 11204 23044
rect 11152 23001 11161 23035
rect 11161 23001 11195 23035
rect 11195 23001 11204 23035
rect 11152 22992 11204 23001
rect 4896 22967 4948 22976
rect 4896 22933 4905 22967
rect 4905 22933 4939 22967
rect 4939 22933 4948 22967
rect 4896 22924 4948 22933
rect 6368 22967 6420 22976
rect 6368 22933 6377 22967
rect 6377 22933 6411 22967
rect 6411 22933 6420 22967
rect 6368 22924 6420 22933
rect 6644 22924 6696 22976
rect 9036 22924 9088 22976
rect 12072 23060 12124 23112
rect 12348 23060 12400 23112
rect 13084 23128 13136 23180
rect 12532 23060 12584 23112
rect 12716 23103 12768 23112
rect 12716 23069 12725 23103
rect 12725 23069 12759 23103
rect 12759 23069 12768 23103
rect 12716 23060 12768 23069
rect 12992 23060 13044 23112
rect 13820 23128 13872 23180
rect 16488 23171 16540 23180
rect 16488 23137 16497 23171
rect 16497 23137 16531 23171
rect 16531 23137 16540 23171
rect 16488 23128 16540 23137
rect 19156 23264 19208 23316
rect 19616 23264 19668 23316
rect 19708 23196 19760 23248
rect 21088 23307 21140 23316
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 21548 23264 21600 23316
rect 21272 23196 21324 23248
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 13176 22992 13228 23044
rect 15568 23060 15620 23112
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 13360 22924 13412 22976
rect 13728 22924 13780 22976
rect 14556 22924 14608 22976
rect 16580 23060 16632 23112
rect 17776 23060 17828 23112
rect 19156 23128 19208 23180
rect 18972 23060 19024 23112
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 20536 23128 20588 23180
rect 16028 22924 16080 22976
rect 17040 22924 17092 22976
rect 18604 22992 18656 23044
rect 17960 22967 18012 22976
rect 17960 22933 17969 22967
rect 17969 22933 18003 22967
rect 18003 22933 18012 22967
rect 17960 22924 18012 22933
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 20168 23103 20220 23112
rect 20168 23069 20177 23103
rect 20177 23069 20211 23103
rect 20211 23069 20220 23103
rect 20996 23128 21048 23180
rect 20168 23060 20220 23069
rect 21180 23060 21232 23112
rect 21272 23060 21324 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 22192 23196 22244 23248
rect 20260 22992 20312 23044
rect 20628 22992 20680 23044
rect 20812 23035 20864 23044
rect 20812 23001 20821 23035
rect 20821 23001 20855 23035
rect 20855 23001 20864 23035
rect 20812 22992 20864 23001
rect 21732 22992 21784 23044
rect 25228 23103 25280 23112
rect 25228 23069 25237 23103
rect 25237 23069 25271 23103
rect 25271 23069 25280 23103
rect 25228 23060 25280 23069
rect 25872 23103 25924 23112
rect 25872 23069 25881 23103
rect 25881 23069 25915 23103
rect 25915 23069 25924 23103
rect 25872 23060 25924 23069
rect 21180 22967 21232 22976
rect 21180 22933 21189 22967
rect 21189 22933 21223 22967
rect 21223 22933 21232 22967
rect 21180 22924 21232 22933
rect 21916 22967 21968 22976
rect 21916 22933 21925 22967
rect 21925 22933 21959 22967
rect 21959 22933 21968 22967
rect 21916 22924 21968 22933
rect 25596 22924 25648 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 2504 22763 2556 22772
rect 2504 22729 2513 22763
rect 2513 22729 2547 22763
rect 2547 22729 2556 22763
rect 2504 22720 2556 22729
rect 2596 22720 2648 22772
rect 4988 22720 5040 22772
rect 5264 22720 5316 22772
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 3148 22559 3200 22568
rect 3148 22525 3157 22559
rect 3157 22525 3191 22559
rect 3191 22525 3200 22559
rect 3148 22516 3200 22525
rect 3608 22627 3660 22636
rect 3608 22593 3617 22627
rect 3617 22593 3651 22627
rect 3651 22593 3660 22627
rect 3608 22584 3660 22593
rect 4804 22652 4856 22704
rect 6644 22652 6696 22704
rect 7012 22763 7064 22772
rect 7012 22729 7021 22763
rect 7021 22729 7055 22763
rect 7055 22729 7064 22763
rect 7012 22720 7064 22729
rect 7932 22652 7984 22704
rect 11612 22720 11664 22772
rect 13176 22720 13228 22772
rect 14740 22720 14792 22772
rect 16212 22720 16264 22772
rect 8668 22652 8720 22704
rect 12440 22652 12492 22704
rect 13912 22652 13964 22704
rect 18052 22720 18104 22772
rect 7840 22584 7892 22636
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 3792 22516 3844 22568
rect 4620 22559 4672 22568
rect 4620 22525 4629 22559
rect 4629 22525 4663 22559
rect 4663 22525 4672 22559
rect 4620 22516 4672 22525
rect 6828 22516 6880 22568
rect 7748 22516 7800 22568
rect 11060 22516 11112 22568
rect 1952 22448 2004 22500
rect 8760 22491 8812 22500
rect 8760 22457 8769 22491
rect 8769 22457 8803 22491
rect 8803 22457 8812 22491
rect 8760 22448 8812 22457
rect 11428 22516 11480 22568
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 16028 22627 16080 22636
rect 16028 22593 16037 22627
rect 16037 22593 16071 22627
rect 16071 22593 16080 22627
rect 16028 22584 16080 22593
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 17224 22695 17276 22704
rect 17224 22661 17258 22695
rect 17258 22661 17276 22695
rect 17224 22652 17276 22661
rect 17960 22652 18012 22704
rect 18604 22652 18656 22704
rect 18328 22627 18380 22636
rect 12072 22516 12124 22568
rect 15568 22516 15620 22568
rect 16672 22516 16724 22568
rect 12256 22448 12308 22500
rect 3608 22380 3660 22432
rect 4620 22380 4672 22432
rect 4896 22380 4948 22432
rect 5356 22380 5408 22432
rect 11704 22380 11756 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 11980 22380 12032 22432
rect 13820 22380 13872 22432
rect 15476 22380 15528 22432
rect 17040 22559 17092 22568
rect 17040 22525 17049 22559
rect 17049 22525 17083 22559
rect 17083 22525 17092 22559
rect 17040 22516 17092 22525
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 18328 22584 18380 22593
rect 17592 22516 17644 22568
rect 18696 22627 18748 22636
rect 18696 22593 18705 22627
rect 18705 22593 18739 22627
rect 18739 22593 18748 22627
rect 18696 22584 18748 22593
rect 18972 22627 19024 22636
rect 18972 22593 18981 22627
rect 18981 22593 19015 22627
rect 19015 22593 19024 22627
rect 18972 22584 19024 22593
rect 19156 22584 19208 22636
rect 19340 22627 19392 22636
rect 19340 22593 19349 22627
rect 19349 22593 19383 22627
rect 19383 22593 19392 22627
rect 19340 22584 19392 22593
rect 19616 22652 19668 22704
rect 20812 22720 20864 22772
rect 21916 22720 21968 22772
rect 20352 22652 20404 22704
rect 20812 22584 20864 22636
rect 23480 22584 23532 22636
rect 24400 22584 24452 22636
rect 25228 22584 25280 22636
rect 25596 22627 25648 22636
rect 25596 22593 25605 22627
rect 25605 22593 25639 22627
rect 25639 22593 25648 22627
rect 25596 22584 25648 22593
rect 17684 22448 17736 22500
rect 19432 22516 19484 22568
rect 21640 22516 21692 22568
rect 24768 22516 24820 22568
rect 17868 22423 17920 22432
rect 17868 22389 17877 22423
rect 17877 22389 17911 22423
rect 17911 22389 17920 22423
rect 17868 22380 17920 22389
rect 20352 22448 20404 22500
rect 21088 22448 21140 22500
rect 19156 22423 19208 22432
rect 19156 22389 19165 22423
rect 19165 22389 19199 22423
rect 19199 22389 19208 22423
rect 19156 22380 19208 22389
rect 19524 22380 19576 22432
rect 19800 22423 19852 22432
rect 19800 22389 19809 22423
rect 19809 22389 19843 22423
rect 19843 22389 19852 22423
rect 19800 22380 19852 22389
rect 19984 22423 20036 22432
rect 19984 22389 19993 22423
rect 19993 22389 20027 22423
rect 20027 22389 20036 22423
rect 19984 22380 20036 22389
rect 20720 22380 20772 22432
rect 20996 22380 21048 22432
rect 21180 22380 21232 22432
rect 21364 22380 21416 22432
rect 21456 22423 21508 22432
rect 21456 22389 21465 22423
rect 21465 22389 21499 22423
rect 21499 22389 21508 22423
rect 21456 22380 21508 22389
rect 25780 22423 25832 22432
rect 25780 22389 25789 22423
rect 25789 22389 25823 22423
rect 25823 22389 25832 22423
rect 25780 22380 25832 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 3608 22176 3660 22228
rect 4528 22176 4580 22228
rect 4712 22176 4764 22228
rect 5448 22176 5500 22228
rect 2780 22108 2832 22160
rect 3700 22108 3752 22160
rect 3792 22108 3844 22160
rect 5172 22108 5224 22160
rect 6368 22108 6420 22160
rect 17868 22176 17920 22228
rect 18972 22176 19024 22228
rect 19340 22176 19392 22228
rect 19616 22176 19668 22228
rect 20168 22176 20220 22228
rect 2504 22083 2556 22092
rect 2504 22049 2513 22083
rect 2513 22049 2547 22083
rect 2547 22049 2556 22083
rect 2504 22040 2556 22049
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 2412 21972 2464 21981
rect 2688 21972 2740 22024
rect 3148 21972 3200 22024
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 3608 21904 3660 21956
rect 2136 21879 2188 21888
rect 2136 21845 2145 21879
rect 2145 21845 2179 21879
rect 2179 21845 2188 21879
rect 2136 21836 2188 21845
rect 4896 22015 4948 22024
rect 4896 21981 4905 22015
rect 4905 21981 4939 22015
rect 4939 21981 4948 22015
rect 4896 21972 4948 21981
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 8668 22108 8720 22160
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 12256 22108 12308 22160
rect 17316 22108 17368 22160
rect 19432 22108 19484 22160
rect 11152 22040 11204 22092
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 7104 21972 7156 22024
rect 9128 21972 9180 22024
rect 5356 21836 5408 21888
rect 5908 21836 5960 21888
rect 6828 21836 6880 21888
rect 7840 21879 7892 21888
rect 7840 21845 7849 21879
rect 7849 21845 7883 21879
rect 7883 21845 7892 21879
rect 7840 21836 7892 21845
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 8208 21836 8260 21845
rect 10140 21836 10192 21888
rect 11244 21972 11296 22024
rect 11428 22015 11480 22024
rect 11428 21981 11437 22015
rect 11437 21981 11471 22015
rect 11471 21981 11480 22015
rect 11428 21972 11480 21981
rect 11704 21904 11756 21956
rect 11888 21972 11940 22024
rect 16120 22040 16172 22092
rect 16672 22040 16724 22092
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 13544 21972 13596 22024
rect 15568 21972 15620 22024
rect 17040 21972 17092 22024
rect 16764 21904 16816 21956
rect 17224 21972 17276 22024
rect 17592 21972 17644 22024
rect 18052 22040 18104 22092
rect 20352 22083 20404 22092
rect 19064 21972 19116 22024
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 20720 22108 20772 22160
rect 21364 22176 21416 22228
rect 21548 22219 21600 22228
rect 21548 22185 21557 22219
rect 21557 22185 21591 22219
rect 21591 22185 21600 22219
rect 21548 22176 21600 22185
rect 21916 22176 21968 22228
rect 21180 22108 21232 22160
rect 21272 22040 21324 22092
rect 22100 22040 22152 22092
rect 24400 22219 24452 22228
rect 24400 22185 24409 22219
rect 24409 22185 24443 22219
rect 24443 22185 24452 22219
rect 24400 22176 24452 22185
rect 22744 22040 22796 22092
rect 23480 22040 23532 22092
rect 19708 21904 19760 21956
rect 20628 21972 20680 22024
rect 20812 21972 20864 22024
rect 11152 21836 11204 21888
rect 11888 21836 11940 21888
rect 13176 21836 13228 21888
rect 14464 21836 14516 21888
rect 14648 21836 14700 21888
rect 17224 21836 17276 21888
rect 19800 21836 19852 21888
rect 19892 21879 19944 21888
rect 19892 21845 19901 21879
rect 19901 21845 19935 21879
rect 19935 21845 19944 21879
rect 19892 21836 19944 21845
rect 20812 21879 20864 21888
rect 20812 21845 20821 21879
rect 20821 21845 20855 21879
rect 20855 21845 20864 21879
rect 20812 21836 20864 21845
rect 21364 21904 21416 21956
rect 21548 21950 21600 22002
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 21180 21836 21232 21888
rect 23664 21904 23716 21956
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 22008 21836 22060 21888
rect 22376 21836 22428 21888
rect 23940 21836 23992 21888
rect 25412 21879 25464 21888
rect 25412 21845 25421 21879
rect 25421 21845 25455 21879
rect 25455 21845 25464 21879
rect 25412 21836 25464 21845
rect 25964 21836 26016 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 3608 21675 3660 21684
rect 3608 21641 3617 21675
rect 3617 21641 3651 21675
rect 3651 21641 3660 21675
rect 3608 21632 3660 21641
rect 2136 21564 2188 21616
rect 848 21496 900 21548
rect 3332 21496 3384 21548
rect 3792 21496 3844 21548
rect 6920 21632 6972 21684
rect 9128 21632 9180 21684
rect 11796 21632 11848 21684
rect 11888 21675 11940 21684
rect 11888 21641 11897 21675
rect 11897 21641 11931 21675
rect 11931 21641 11940 21675
rect 11888 21632 11940 21641
rect 12256 21632 12308 21684
rect 12808 21632 12860 21684
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 1952 21428 2004 21480
rect 6736 21428 6788 21480
rect 3240 21292 3292 21344
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 3424 21292 3476 21301
rect 6460 21292 6512 21344
rect 6644 21292 6696 21344
rect 7012 21496 7064 21548
rect 8300 21564 8352 21616
rect 12716 21564 12768 21616
rect 13452 21564 13504 21616
rect 7104 21403 7156 21412
rect 7104 21369 7113 21403
rect 7113 21369 7147 21403
rect 7147 21369 7156 21403
rect 7104 21360 7156 21369
rect 8208 21496 8260 21548
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 12900 21496 12952 21548
rect 9588 21428 9640 21480
rect 9496 21292 9548 21344
rect 12256 21292 12308 21344
rect 14832 21496 14884 21548
rect 15660 21496 15712 21548
rect 19984 21496 20036 21548
rect 22192 21632 22244 21684
rect 23388 21632 23440 21684
rect 20996 21564 21048 21616
rect 22284 21564 22336 21616
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 21180 21496 21232 21548
rect 21272 21496 21324 21548
rect 21732 21496 21784 21548
rect 21916 21496 21968 21548
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 19892 21471 19944 21480
rect 19892 21437 19901 21471
rect 19901 21437 19935 21471
rect 19935 21437 19944 21471
rect 19892 21428 19944 21437
rect 20352 21428 20404 21480
rect 20720 21428 20772 21480
rect 19984 21403 20036 21412
rect 19984 21369 19993 21403
rect 19993 21369 20027 21403
rect 20027 21369 20036 21403
rect 19984 21360 20036 21369
rect 13636 21292 13688 21344
rect 13820 21292 13872 21344
rect 19156 21292 19208 21344
rect 21180 21360 21232 21412
rect 21640 21428 21692 21480
rect 20168 21292 20220 21344
rect 20812 21292 20864 21344
rect 21088 21292 21140 21344
rect 21272 21335 21324 21344
rect 21272 21301 21281 21335
rect 21281 21301 21315 21335
rect 21315 21301 21324 21335
rect 21272 21292 21324 21301
rect 21824 21360 21876 21412
rect 23204 21496 23256 21548
rect 23572 21496 23624 21548
rect 23756 21539 23808 21548
rect 23756 21505 23765 21539
rect 23765 21505 23799 21539
rect 23799 21505 23808 21539
rect 23756 21496 23808 21505
rect 24032 21539 24084 21548
rect 24032 21505 24066 21539
rect 24066 21505 24084 21539
rect 24032 21496 24084 21505
rect 22928 21471 22980 21480
rect 22928 21437 22937 21471
rect 22937 21437 22971 21471
rect 22971 21437 22980 21471
rect 22928 21428 22980 21437
rect 23664 21403 23716 21412
rect 23664 21369 23673 21403
rect 23673 21369 23707 21403
rect 23707 21369 23716 21403
rect 23664 21360 23716 21369
rect 22560 21292 22612 21344
rect 25228 21335 25280 21344
rect 25228 21301 25237 21335
rect 25237 21301 25271 21335
rect 25271 21301 25280 21335
rect 25228 21292 25280 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 3240 20952 3292 21004
rect 5356 21088 5408 21140
rect 11244 21131 11296 21140
rect 11244 21097 11253 21131
rect 11253 21097 11287 21131
rect 11287 21097 11296 21131
rect 11244 21088 11296 21097
rect 11980 21088 12032 21140
rect 12716 21088 12768 21140
rect 12808 21088 12860 21140
rect 13452 21088 13504 21140
rect 14096 21088 14148 21140
rect 14832 21088 14884 21140
rect 19984 21088 20036 21140
rect 5724 21020 5776 21072
rect 5816 21020 5868 21072
rect 6644 21020 6696 21072
rect 1952 20884 2004 20936
rect 2412 20884 2464 20936
rect 2872 20884 2924 20936
rect 3424 20884 3476 20936
rect 4068 20884 4120 20936
rect 6368 20952 6420 21004
rect 6460 20952 6512 21004
rect 2136 20859 2188 20868
rect 2136 20825 2170 20859
rect 2170 20825 2188 20859
rect 2136 20816 2188 20825
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 4804 20816 4856 20868
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6000 20884 6052 20936
rect 6552 20884 6604 20936
rect 9496 21063 9548 21072
rect 9496 21029 9505 21063
rect 9505 21029 9539 21063
rect 9539 21029 9548 21063
rect 9496 21020 9548 21029
rect 12624 21063 12676 21072
rect 12624 21029 12633 21063
rect 12633 21029 12667 21063
rect 12667 21029 12676 21063
rect 12624 21020 12676 21029
rect 14372 21020 14424 21072
rect 9588 20884 9640 20936
rect 10140 20927 10192 20936
rect 10140 20893 10174 20927
rect 10174 20893 10192 20927
rect 10140 20884 10192 20893
rect 12716 20952 12768 21004
rect 12992 20995 13044 21004
rect 12992 20961 13001 20995
rect 13001 20961 13035 20995
rect 13035 20961 13044 20995
rect 12992 20952 13044 20961
rect 13452 20952 13504 21004
rect 13636 20995 13688 21004
rect 13636 20961 13645 20995
rect 13645 20961 13679 20995
rect 13679 20961 13688 20995
rect 13636 20952 13688 20961
rect 14280 20995 14332 21004
rect 14280 20961 14289 20995
rect 14289 20961 14323 20995
rect 14323 20961 14332 20995
rect 14280 20952 14332 20961
rect 14464 20995 14516 21004
rect 14464 20961 14473 20995
rect 14473 20961 14507 20995
rect 14507 20961 14516 20995
rect 14464 20952 14516 20961
rect 12164 20884 12216 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 12808 20929 12860 20936
rect 12808 20895 12817 20929
rect 12817 20895 12851 20929
rect 12851 20895 12860 20929
rect 12808 20884 12860 20895
rect 6736 20816 6788 20868
rect 4620 20791 4672 20800
rect 4620 20757 4629 20791
rect 4629 20757 4663 20791
rect 4663 20757 4672 20791
rect 4620 20748 4672 20757
rect 5632 20791 5684 20800
rect 5632 20757 5641 20791
rect 5641 20757 5675 20791
rect 5675 20757 5684 20791
rect 5632 20748 5684 20757
rect 6828 20791 6880 20800
rect 6828 20757 6837 20791
rect 6837 20757 6871 20791
rect 6871 20757 6880 20791
rect 6828 20748 6880 20757
rect 7380 20791 7432 20800
rect 7380 20757 7389 20791
rect 7389 20757 7423 20791
rect 7423 20757 7432 20791
rect 7380 20748 7432 20757
rect 8300 20816 8352 20868
rect 8392 20816 8444 20868
rect 8944 20859 8996 20868
rect 8944 20825 8953 20859
rect 8953 20825 8987 20859
rect 8987 20825 8996 20859
rect 8944 20816 8996 20825
rect 9036 20816 9088 20868
rect 9312 20791 9364 20800
rect 9312 20757 9321 20791
rect 9321 20757 9355 20791
rect 9355 20757 9364 20791
rect 9312 20748 9364 20757
rect 11520 20791 11572 20800
rect 11520 20757 11529 20791
rect 11529 20757 11563 20791
rect 11563 20757 11572 20791
rect 11520 20748 11572 20757
rect 11888 20791 11940 20800
rect 11888 20757 11897 20791
rect 11897 20757 11931 20791
rect 11931 20757 11940 20791
rect 11888 20748 11940 20757
rect 13728 20884 13780 20936
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 17408 20952 17460 21004
rect 19064 20952 19116 21004
rect 20720 21131 20772 21140
rect 20720 21097 20729 21131
rect 20729 21097 20763 21131
rect 20763 21097 20772 21131
rect 20720 21088 20772 21097
rect 20628 21020 20680 21072
rect 21180 21088 21232 21140
rect 22284 21088 22336 21140
rect 23940 21088 23992 21140
rect 24032 21088 24084 21140
rect 17316 20884 17368 20936
rect 17500 20884 17552 20936
rect 19156 20816 19208 20868
rect 19708 20927 19760 20936
rect 19708 20893 19717 20927
rect 19717 20893 19751 20927
rect 19751 20893 19760 20927
rect 19708 20884 19760 20893
rect 19892 20927 19944 20936
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 20628 20884 20680 20936
rect 21364 21020 21416 21072
rect 21640 21020 21692 21072
rect 23756 20952 23808 21004
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 21272 20884 21324 20936
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 21732 20884 21784 20936
rect 22928 20884 22980 20936
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 25228 20884 25280 20936
rect 20720 20816 20772 20868
rect 15200 20748 15252 20800
rect 16672 20791 16724 20800
rect 16672 20757 16681 20791
rect 16681 20757 16715 20791
rect 16715 20757 16724 20791
rect 16672 20748 16724 20757
rect 18696 20748 18748 20800
rect 19432 20748 19484 20800
rect 19800 20791 19852 20800
rect 19800 20757 19809 20791
rect 19809 20757 19843 20791
rect 19843 20757 19852 20791
rect 21548 20816 21600 20868
rect 22284 20859 22336 20868
rect 22284 20825 22293 20859
rect 22293 20825 22327 20859
rect 22327 20825 22336 20859
rect 22284 20816 22336 20825
rect 22560 20816 22612 20868
rect 24676 20859 24728 20868
rect 24676 20825 24710 20859
rect 24710 20825 24728 20859
rect 19800 20748 19852 20757
rect 22008 20791 22060 20800
rect 22008 20757 22017 20791
rect 22017 20757 22051 20791
rect 22051 20757 22060 20791
rect 22008 20748 22060 20757
rect 22652 20748 22704 20800
rect 24676 20816 24728 20825
rect 23664 20748 23716 20800
rect 25780 20791 25832 20800
rect 25780 20757 25789 20791
rect 25789 20757 25823 20791
rect 25823 20757 25832 20791
rect 25780 20748 25832 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 2136 20544 2188 20596
rect 2320 20587 2372 20596
rect 2320 20553 2329 20587
rect 2329 20553 2363 20587
rect 2363 20553 2372 20587
rect 2320 20544 2372 20553
rect 2412 20544 2464 20596
rect 2780 20476 2832 20528
rect 3240 20476 3292 20528
rect 3792 20519 3844 20528
rect 3792 20485 3801 20519
rect 3801 20485 3835 20519
rect 3835 20485 3844 20519
rect 3792 20476 3844 20485
rect 4068 20476 4120 20528
rect 7380 20544 7432 20596
rect 9312 20544 9364 20596
rect 1952 20451 2004 20460
rect 1952 20417 1961 20451
rect 1961 20417 1995 20451
rect 1995 20417 2004 20451
rect 1952 20408 2004 20417
rect 2504 20408 2556 20460
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 3424 20340 3476 20392
rect 2872 20272 2924 20324
rect 2228 20204 2280 20256
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 4528 20408 4580 20460
rect 4620 20451 4672 20460
rect 4620 20417 4629 20451
rect 4629 20417 4663 20451
rect 4663 20417 4672 20451
rect 4620 20408 4672 20417
rect 4712 20451 4764 20460
rect 4712 20417 4721 20451
rect 4721 20417 4755 20451
rect 4755 20417 4764 20451
rect 4712 20408 4764 20417
rect 8300 20476 8352 20528
rect 9036 20476 9088 20528
rect 9128 20476 9180 20528
rect 12532 20544 12584 20596
rect 12440 20476 12492 20528
rect 12624 20519 12676 20528
rect 12624 20485 12642 20519
rect 12642 20485 12676 20519
rect 12900 20544 12952 20596
rect 13820 20544 13872 20596
rect 14004 20587 14056 20596
rect 14004 20553 14013 20587
rect 14013 20553 14047 20587
rect 14047 20553 14056 20587
rect 14004 20544 14056 20553
rect 15200 20587 15252 20596
rect 15200 20553 15209 20587
rect 15209 20553 15243 20587
rect 15243 20553 15252 20587
rect 15200 20544 15252 20553
rect 17408 20544 17460 20596
rect 12624 20476 12676 20485
rect 14096 20476 14148 20528
rect 5080 20340 5132 20392
rect 10508 20340 10560 20392
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 13544 20408 13596 20460
rect 15016 20476 15068 20528
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 15384 20408 15436 20460
rect 14464 20383 14516 20392
rect 14464 20349 14473 20383
rect 14473 20349 14507 20383
rect 14507 20349 14516 20383
rect 14464 20340 14516 20349
rect 17316 20408 17368 20460
rect 19800 20544 19852 20596
rect 20628 20544 20680 20596
rect 21364 20587 21416 20596
rect 21364 20553 21373 20587
rect 21373 20553 21407 20587
rect 21407 20553 21416 20587
rect 21364 20544 21416 20553
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 19432 20476 19484 20528
rect 5172 20204 5224 20256
rect 8668 20204 8720 20256
rect 12532 20204 12584 20256
rect 13360 20272 13412 20324
rect 15292 20272 15344 20324
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 19708 20408 19760 20460
rect 20168 20408 20220 20460
rect 19892 20340 19944 20392
rect 19800 20272 19852 20324
rect 20536 20272 20588 20324
rect 20720 20340 20772 20392
rect 22192 20476 22244 20528
rect 22928 20544 22980 20596
rect 23112 20544 23164 20596
rect 23664 20544 23716 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 25596 20544 25648 20596
rect 21640 20408 21692 20460
rect 21916 20408 21968 20460
rect 21088 20340 21140 20392
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 22192 20383 22244 20392
rect 22192 20349 22201 20383
rect 22201 20349 22235 20383
rect 22235 20349 22244 20383
rect 22192 20340 22244 20349
rect 12992 20204 13044 20256
rect 13452 20204 13504 20256
rect 14280 20204 14332 20256
rect 15200 20204 15252 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20352 20204 20404 20213
rect 21272 20272 21324 20324
rect 22008 20272 22060 20324
rect 22468 20408 22520 20460
rect 23112 20408 23164 20460
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23572 20451 23624 20460
rect 23572 20417 23581 20451
rect 23581 20417 23615 20451
rect 23615 20417 23624 20451
rect 23572 20408 23624 20417
rect 25780 20408 25832 20460
rect 22836 20340 22888 20392
rect 23112 20204 23164 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 1952 20000 2004 20052
rect 3240 20000 3292 20052
rect 3792 20000 3844 20052
rect 6828 20000 6880 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 14464 20000 14516 20052
rect 17132 20000 17184 20052
rect 17500 20000 17552 20052
rect 19432 20000 19484 20052
rect 3608 19864 3660 19916
rect 4068 19864 4120 19916
rect 2780 19796 2832 19848
rect 3240 19796 3292 19848
rect 3884 19796 3936 19848
rect 4620 19796 4672 19848
rect 5080 19839 5132 19848
rect 5080 19805 5089 19839
rect 5089 19805 5123 19839
rect 5123 19805 5132 19839
rect 5080 19796 5132 19805
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 5632 19796 5684 19848
rect 5724 19796 5776 19848
rect 7748 19907 7800 19916
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 8300 19932 8352 19984
rect 8484 19932 8536 19984
rect 19340 19932 19392 19984
rect 8944 19864 8996 19916
rect 15660 19907 15712 19916
rect 15660 19873 15669 19907
rect 15669 19873 15703 19907
rect 15703 19873 15712 19907
rect 15660 19864 15712 19873
rect 19064 19864 19116 19916
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 11060 19796 11112 19848
rect 11520 19796 11572 19848
rect 12072 19796 12124 19848
rect 12900 19796 12952 19848
rect 6828 19728 6880 19780
rect 11428 19728 11480 19780
rect 11888 19728 11940 19780
rect 14096 19796 14148 19848
rect 16672 19796 16724 19848
rect 18052 19796 18104 19848
rect 19248 19839 19300 19848
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 19892 19796 19944 19848
rect 20812 20000 20864 20052
rect 21916 20000 21968 20052
rect 22192 20043 22244 20052
rect 22192 20009 22201 20043
rect 22201 20009 22235 20043
rect 22235 20009 22244 20043
rect 22192 20000 22244 20009
rect 20996 19932 21048 19984
rect 21364 19932 21416 19984
rect 21180 19864 21232 19916
rect 20996 19839 21048 19848
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 14832 19728 14884 19780
rect 2228 19660 2280 19712
rect 5632 19660 5684 19712
rect 5816 19703 5868 19712
rect 5816 19669 5825 19703
rect 5825 19669 5859 19703
rect 5859 19669 5868 19703
rect 5816 19660 5868 19669
rect 5908 19703 5960 19712
rect 5908 19669 5917 19703
rect 5917 19669 5951 19703
rect 5951 19669 5960 19703
rect 5908 19660 5960 19669
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 8668 19660 8720 19712
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 18328 19660 18380 19712
rect 19248 19660 19300 19712
rect 21364 19796 21416 19848
rect 21640 19839 21692 19848
rect 21640 19805 21649 19839
rect 21649 19805 21683 19839
rect 21683 19805 21692 19839
rect 21640 19796 21692 19805
rect 23296 19932 23348 19984
rect 22468 19864 22520 19916
rect 22100 19796 22152 19848
rect 22284 19796 22336 19848
rect 22560 19839 22612 19848
rect 22560 19805 22569 19839
rect 22569 19805 22603 19839
rect 22603 19805 22612 19839
rect 22560 19796 22612 19805
rect 23940 19839 23992 19848
rect 23940 19805 23949 19839
rect 23949 19805 23983 19839
rect 23983 19805 23992 19839
rect 23940 19796 23992 19805
rect 25320 19796 25372 19848
rect 22376 19771 22428 19780
rect 22376 19737 22385 19771
rect 22385 19737 22419 19771
rect 22419 19737 22428 19771
rect 22376 19728 22428 19737
rect 21272 19660 21324 19712
rect 21824 19660 21876 19712
rect 23572 19660 23624 19712
rect 23848 19660 23900 19712
rect 24124 19703 24176 19712
rect 24124 19669 24133 19703
rect 24133 19669 24167 19703
rect 24167 19669 24176 19703
rect 24124 19660 24176 19669
rect 24400 19703 24452 19712
rect 24400 19669 24409 19703
rect 24409 19669 24443 19703
rect 24443 19669 24452 19703
rect 24400 19660 24452 19669
rect 24492 19660 24544 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 12440 19456 12492 19508
rect 13912 19499 13964 19508
rect 13912 19465 13921 19499
rect 13921 19465 13955 19499
rect 13955 19465 13964 19499
rect 13912 19456 13964 19465
rect 14464 19456 14516 19508
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 20996 19456 21048 19508
rect 2320 19388 2372 19440
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 3148 19388 3200 19440
rect 3792 19363 3844 19372
rect 3792 19329 3801 19363
rect 3801 19329 3835 19363
rect 3835 19329 3844 19363
rect 3792 19320 3844 19329
rect 4068 19320 4120 19372
rect 4712 19320 4764 19372
rect 2780 19252 2832 19304
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 4620 19252 4672 19304
rect 5816 19388 5868 19440
rect 5908 19320 5960 19372
rect 6000 19320 6052 19372
rect 7840 19388 7892 19440
rect 8208 19388 8260 19440
rect 6552 19320 6604 19372
rect 6920 19320 6972 19372
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 11428 19320 11480 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 14096 19320 14148 19372
rect 16672 19320 16724 19372
rect 17224 19363 17276 19372
rect 17224 19329 17233 19363
rect 17233 19329 17267 19363
rect 17267 19329 17276 19363
rect 17224 19320 17276 19329
rect 19432 19388 19484 19440
rect 22192 19456 22244 19508
rect 22468 19499 22520 19508
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 23940 19456 23992 19508
rect 21640 19388 21692 19440
rect 25320 19456 25372 19508
rect 25780 19499 25832 19508
rect 25780 19465 25789 19499
rect 25789 19465 25823 19499
rect 25823 19465 25832 19499
rect 25780 19456 25832 19465
rect 19248 19320 19300 19372
rect 21916 19320 21968 19372
rect 24400 19388 24452 19440
rect 24860 19388 24912 19440
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 8668 19252 8720 19304
rect 7472 19184 7524 19236
rect 7932 19184 7984 19236
rect 8116 19184 8168 19236
rect 10416 19184 10468 19236
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 4804 19116 4856 19168
rect 6000 19116 6052 19168
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 10324 19116 10376 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 13268 19295 13320 19304
rect 13268 19261 13277 19295
rect 13277 19261 13311 19295
rect 13311 19261 13320 19295
rect 13268 19252 13320 19261
rect 13636 19252 13688 19304
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 15660 19252 15712 19304
rect 18052 19252 18104 19304
rect 13820 19184 13872 19236
rect 22100 19184 22152 19236
rect 14004 19159 14056 19168
rect 14004 19125 14013 19159
rect 14013 19125 14047 19159
rect 14047 19125 14056 19159
rect 14004 19116 14056 19125
rect 21088 19159 21140 19168
rect 21088 19125 21097 19159
rect 21097 19125 21131 19159
rect 21131 19125 21140 19159
rect 21088 19116 21140 19125
rect 21180 19116 21232 19168
rect 21548 19116 21600 19168
rect 22008 19116 22060 19168
rect 23756 19320 23808 19372
rect 25504 19363 25556 19372
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 22560 19116 22612 19168
rect 25320 19159 25372 19168
rect 25320 19125 25329 19159
rect 25329 19125 25363 19159
rect 25363 19125 25372 19159
rect 25320 19116 25372 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 4160 18912 4212 18964
rect 5080 18912 5132 18964
rect 2688 18887 2740 18896
rect 2688 18853 2697 18887
rect 2697 18853 2731 18887
rect 2731 18853 2740 18887
rect 10508 18912 10560 18964
rect 12532 18912 12584 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 22468 18912 22520 18964
rect 24492 18912 24544 18964
rect 2688 18844 2740 18853
rect 2504 18776 2556 18828
rect 2596 18776 2648 18828
rect 3148 18819 3200 18828
rect 3148 18785 3157 18819
rect 3157 18785 3191 18819
rect 3191 18785 3200 18819
rect 3148 18776 3200 18785
rect 7840 18844 7892 18896
rect 8484 18844 8536 18896
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 5724 18776 5776 18828
rect 848 18708 900 18760
rect 2320 18708 2372 18760
rect 3792 18708 3844 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 2780 18640 2832 18692
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 5356 18751 5408 18760
rect 5356 18717 5387 18751
rect 5387 18717 5408 18751
rect 5356 18708 5408 18717
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 5540 18640 5592 18692
rect 6552 18708 6604 18760
rect 6736 18776 6788 18828
rect 7380 18708 7432 18760
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 10784 18844 10836 18896
rect 12440 18844 12492 18896
rect 12348 18776 12400 18828
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 4436 18572 4488 18624
rect 6460 18683 6512 18692
rect 6460 18649 6469 18683
rect 6469 18649 6503 18683
rect 6503 18649 6512 18683
rect 6460 18640 6512 18649
rect 8944 18708 8996 18760
rect 10232 18708 10284 18760
rect 13084 18708 13136 18760
rect 22560 18844 22612 18896
rect 13360 18776 13412 18828
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 22008 18776 22060 18828
rect 5908 18572 5960 18624
rect 6276 18615 6328 18624
rect 6276 18581 6285 18615
rect 6285 18581 6319 18615
rect 6319 18581 6328 18615
rect 6276 18572 6328 18581
rect 7564 18615 7616 18624
rect 7564 18581 7573 18615
rect 7573 18581 7607 18615
rect 7607 18581 7616 18615
rect 7564 18572 7616 18581
rect 8392 18572 8444 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 9680 18640 9732 18692
rect 12072 18683 12124 18692
rect 12072 18649 12081 18683
rect 12081 18649 12115 18683
rect 12115 18649 12124 18683
rect 12072 18640 12124 18649
rect 12256 18683 12308 18692
rect 12256 18649 12281 18683
rect 12281 18649 12308 18683
rect 13636 18708 13688 18760
rect 14464 18708 14516 18760
rect 14556 18708 14608 18760
rect 16856 18708 16908 18760
rect 20720 18708 20772 18760
rect 21456 18708 21508 18760
rect 21548 18708 21600 18760
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 23572 18776 23624 18828
rect 12256 18640 12308 18649
rect 11704 18615 11756 18624
rect 11704 18581 11729 18615
rect 11729 18581 11756 18615
rect 11704 18572 11756 18581
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 17868 18640 17920 18692
rect 12992 18572 13044 18624
rect 15568 18572 15620 18624
rect 16028 18572 16080 18624
rect 17132 18572 17184 18624
rect 18604 18572 18656 18624
rect 19616 18572 19668 18624
rect 20260 18572 20312 18624
rect 21364 18572 21416 18624
rect 21640 18615 21692 18624
rect 21640 18581 21649 18615
rect 21649 18581 21683 18615
rect 21683 18581 21692 18615
rect 21640 18572 21692 18581
rect 21824 18572 21876 18624
rect 22192 18683 22244 18692
rect 22192 18649 22201 18683
rect 22201 18649 22235 18683
rect 22235 18649 22244 18683
rect 22192 18640 22244 18649
rect 22008 18572 22060 18624
rect 23204 18708 23256 18760
rect 23664 18708 23716 18760
rect 25136 18708 25188 18760
rect 25504 18708 25556 18760
rect 22928 18640 22980 18692
rect 24216 18640 24268 18692
rect 24308 18572 24360 18624
rect 24400 18615 24452 18624
rect 24400 18581 24409 18615
rect 24409 18581 24443 18615
rect 24443 18581 24452 18615
rect 24400 18572 24452 18581
rect 24584 18572 24636 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2228 18368 2280 18420
rect 4068 18368 4120 18420
rect 5264 18368 5316 18420
rect 5540 18411 5592 18420
rect 5540 18377 5549 18411
rect 5549 18377 5583 18411
rect 5583 18377 5592 18411
rect 5540 18368 5592 18377
rect 7380 18368 7432 18420
rect 8116 18368 8168 18420
rect 8392 18368 8444 18420
rect 8852 18368 8904 18420
rect 12256 18368 12308 18420
rect 12440 18368 12492 18420
rect 13084 18368 13136 18420
rect 13544 18411 13596 18420
rect 13544 18377 13553 18411
rect 13553 18377 13587 18411
rect 13587 18377 13596 18411
rect 13544 18368 13596 18377
rect 13820 18411 13872 18420
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 19340 18368 19392 18420
rect 20628 18368 20680 18420
rect 21824 18368 21876 18420
rect 23204 18368 23256 18420
rect 25136 18411 25188 18420
rect 25136 18377 25145 18411
rect 25145 18377 25179 18411
rect 25179 18377 25188 18411
rect 25136 18368 25188 18377
rect 25412 18411 25464 18420
rect 25412 18377 25421 18411
rect 25421 18377 25455 18411
rect 25455 18377 25464 18411
rect 25412 18368 25464 18377
rect 2412 18232 2464 18284
rect 2964 18275 3016 18284
rect 2964 18241 2982 18275
rect 2982 18241 3016 18275
rect 2964 18232 3016 18241
rect 3976 18275 4028 18284
rect 3976 18241 3985 18275
rect 3985 18241 4019 18275
rect 4019 18241 4028 18275
rect 3976 18232 4028 18241
rect 4068 18275 4120 18284
rect 4068 18241 4078 18275
rect 4078 18241 4112 18275
rect 4112 18241 4120 18275
rect 4068 18232 4120 18241
rect 4436 18275 4488 18284
rect 4436 18241 4445 18275
rect 4445 18241 4479 18275
rect 4479 18241 4488 18275
rect 4436 18232 4488 18241
rect 5724 18300 5776 18352
rect 6460 18300 6512 18352
rect 7288 18300 7340 18352
rect 5908 18275 5960 18284
rect 5908 18241 5917 18275
rect 5917 18241 5951 18275
rect 5951 18241 5960 18275
rect 5908 18232 5960 18241
rect 6000 18275 6052 18284
rect 6000 18241 6009 18275
rect 6009 18241 6043 18275
rect 6043 18241 6052 18275
rect 6000 18232 6052 18241
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7196 18275 7248 18284
rect 7196 18241 7205 18275
rect 7205 18241 7239 18275
rect 7239 18241 7248 18275
rect 7196 18232 7248 18241
rect 7932 18300 7984 18352
rect 10324 18343 10376 18352
rect 10324 18309 10342 18343
rect 10342 18309 10376 18343
rect 10324 18300 10376 18309
rect 10416 18343 10468 18352
rect 10416 18309 10425 18343
rect 10425 18309 10459 18343
rect 10459 18309 10468 18343
rect 10416 18300 10468 18309
rect 7012 18164 7064 18216
rect 7104 18164 7156 18216
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8576 18232 8628 18284
rect 7748 18164 7800 18216
rect 8208 18207 8260 18216
rect 8208 18173 8217 18207
rect 8217 18173 8251 18207
rect 8251 18173 8260 18207
rect 8208 18164 8260 18173
rect 10140 18164 10192 18216
rect 12256 18232 12308 18284
rect 10508 18164 10560 18216
rect 12348 18164 12400 18216
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13452 18300 13504 18352
rect 15568 18343 15620 18352
rect 15568 18309 15586 18343
rect 15586 18309 15620 18343
rect 15568 18300 15620 18309
rect 13176 18232 13228 18284
rect 14004 18232 14056 18284
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15752 18232 15804 18284
rect 18144 18232 18196 18284
rect 13636 18164 13688 18216
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 19064 18232 19116 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 19892 18232 19944 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 7472 18028 7524 18080
rect 8484 18028 8536 18080
rect 10048 18028 10100 18080
rect 12900 18096 12952 18148
rect 11888 18028 11940 18080
rect 12532 18028 12584 18080
rect 16856 18071 16908 18080
rect 16856 18037 16865 18071
rect 16865 18037 16899 18071
rect 16899 18037 16908 18071
rect 16856 18028 16908 18037
rect 19432 18207 19484 18216
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 19432 18164 19484 18173
rect 20260 18164 20312 18216
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 20076 18096 20128 18148
rect 21456 18232 21508 18284
rect 21640 18275 21692 18284
rect 21640 18241 21649 18275
rect 21649 18241 21683 18275
rect 21683 18241 21692 18275
rect 21640 18232 21692 18241
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 24400 18300 24452 18352
rect 22284 18275 22336 18284
rect 22284 18241 22293 18275
rect 22293 18241 22327 18275
rect 22327 18241 22336 18275
rect 22284 18232 22336 18241
rect 22744 18232 22796 18284
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 25320 18232 25372 18284
rect 25596 18275 25648 18284
rect 25596 18241 25605 18275
rect 25605 18241 25639 18275
rect 25639 18241 25648 18275
rect 25596 18232 25648 18241
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 21916 18096 21968 18148
rect 22744 18096 22796 18148
rect 20444 18028 20496 18080
rect 21272 18028 21324 18080
rect 21640 18028 21692 18080
rect 22100 18028 22152 18080
rect 25780 18071 25832 18080
rect 25780 18037 25789 18071
rect 25789 18037 25823 18071
rect 25823 18037 25832 18071
rect 25780 18028 25832 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2780 17824 2832 17876
rect 3976 17824 4028 17876
rect 5356 17824 5408 17876
rect 6828 17867 6880 17876
rect 4160 17756 4212 17808
rect 6828 17833 6837 17867
rect 6837 17833 6871 17867
rect 6871 17833 6880 17867
rect 6828 17824 6880 17833
rect 6920 17824 6972 17876
rect 9680 17824 9732 17876
rect 12532 17824 12584 17876
rect 12624 17867 12676 17876
rect 12624 17833 12633 17867
rect 12633 17833 12667 17867
rect 12667 17833 12676 17867
rect 12624 17824 12676 17833
rect 13360 17824 13412 17876
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 15200 17824 15252 17876
rect 7196 17756 7248 17808
rect 7748 17756 7800 17808
rect 2320 17620 2372 17672
rect 3976 17620 4028 17672
rect 6276 17688 6328 17740
rect 1952 17552 2004 17604
rect 4160 17595 4212 17604
rect 4160 17561 4169 17595
rect 4169 17561 4203 17595
rect 4203 17561 4212 17595
rect 4160 17552 4212 17561
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 7380 17688 7432 17740
rect 8944 17799 8996 17808
rect 8944 17765 8953 17799
rect 8953 17765 8987 17799
rect 8987 17765 8996 17799
rect 8944 17756 8996 17765
rect 12072 17799 12124 17808
rect 12072 17765 12081 17799
rect 12081 17765 12115 17799
rect 12115 17765 12124 17799
rect 12072 17756 12124 17765
rect 4436 17484 4488 17536
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 8300 17688 8352 17740
rect 8760 17688 8812 17740
rect 7932 17620 7984 17672
rect 10048 17663 10100 17672
rect 10048 17629 10066 17663
rect 10066 17629 10100 17663
rect 10048 17620 10100 17629
rect 10232 17620 10284 17672
rect 8668 17552 8720 17604
rect 10968 17552 11020 17604
rect 11060 17595 11112 17604
rect 11060 17561 11069 17595
rect 11069 17561 11103 17595
rect 11103 17561 11112 17595
rect 11060 17552 11112 17561
rect 17868 17867 17920 17876
rect 17868 17833 17877 17867
rect 17877 17833 17911 17867
rect 17911 17833 17920 17867
rect 17868 17824 17920 17833
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 19800 17867 19852 17876
rect 19800 17833 19809 17867
rect 19809 17833 19843 17867
rect 19843 17833 19852 17867
rect 19800 17824 19852 17833
rect 20536 17824 20588 17876
rect 20996 17824 21048 17876
rect 21272 17824 21324 17876
rect 23572 17824 23624 17876
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 15476 17663 15528 17672
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 16580 17620 16632 17672
rect 17224 17756 17276 17808
rect 22284 17756 22336 17808
rect 18328 17731 18380 17740
rect 18328 17697 18337 17731
rect 18337 17697 18371 17731
rect 18371 17697 18380 17731
rect 18328 17688 18380 17697
rect 17316 17620 17368 17672
rect 17868 17620 17920 17672
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 20904 17688 20956 17740
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 14556 17552 14608 17604
rect 7196 17484 7248 17536
rect 7564 17484 7616 17536
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 7656 17484 7708 17493
rect 12440 17527 12492 17536
rect 12440 17493 12449 17527
rect 12449 17493 12483 17527
rect 12483 17493 12492 17527
rect 12440 17484 12492 17493
rect 17592 17595 17644 17604
rect 17592 17561 17601 17595
rect 17601 17561 17635 17595
rect 17635 17561 17644 17595
rect 17592 17552 17644 17561
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 19708 17484 19760 17536
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 21640 17688 21692 17740
rect 24308 17688 24360 17740
rect 21548 17620 21600 17672
rect 21732 17620 21784 17672
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 23756 17620 23808 17672
rect 25136 17620 25188 17672
rect 21180 17552 21232 17604
rect 21272 17552 21324 17604
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 24032 17484 24084 17536
rect 24492 17484 24544 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3792 17280 3844 17332
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 8576 17280 8628 17332
rect 11060 17280 11112 17332
rect 14740 17280 14792 17332
rect 16580 17280 16632 17332
rect 3792 17144 3844 17196
rect 4436 17187 4488 17196
rect 4436 17153 4449 17187
rect 4449 17153 4488 17187
rect 3884 17076 3936 17128
rect 4436 17144 4488 17153
rect 6276 17144 6328 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 7104 17144 7156 17196
rect 7196 17144 7248 17196
rect 7564 17187 7616 17196
rect 7564 17153 7573 17187
rect 7573 17153 7607 17187
rect 7607 17153 7616 17187
rect 7564 17144 7616 17153
rect 8944 17144 8996 17196
rect 11796 17187 11848 17196
rect 11796 17153 11830 17187
rect 11830 17153 11848 17187
rect 11796 17144 11848 17153
rect 12900 17144 12952 17196
rect 6184 17076 6236 17128
rect 7932 17076 7984 17128
rect 8484 17076 8536 17128
rect 10968 17076 11020 17128
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 16948 17212 17000 17264
rect 17592 17212 17644 17264
rect 18420 17212 18472 17264
rect 19432 17212 19484 17264
rect 15476 17144 15528 17153
rect 5908 17008 5960 17060
rect 6552 16940 6604 16992
rect 6828 16940 6880 16992
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 12256 16940 12308 16992
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 17868 17144 17920 17196
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 18328 17119 18380 17128
rect 18328 17085 18337 17119
rect 18337 17085 18371 17119
rect 18371 17085 18380 17119
rect 18328 17076 18380 17085
rect 21088 17280 21140 17332
rect 21364 17280 21416 17332
rect 22100 17280 22152 17332
rect 22376 17280 22428 17332
rect 25136 17323 25188 17332
rect 25136 17289 25145 17323
rect 25145 17289 25179 17323
rect 25179 17289 25188 17323
rect 25136 17280 25188 17289
rect 25596 17280 25648 17332
rect 19708 17212 19760 17264
rect 20260 17187 20312 17196
rect 20260 17153 20269 17187
rect 20269 17153 20303 17187
rect 20303 17153 20312 17187
rect 20260 17144 20312 17153
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 20720 17144 20772 17196
rect 20904 17144 20956 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 22284 17255 22336 17264
rect 22284 17221 22293 17255
rect 22293 17221 22327 17255
rect 22327 17221 22336 17255
rect 22284 17212 22336 17221
rect 21272 17144 21324 17153
rect 21640 17144 21692 17196
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 18512 17008 18564 17060
rect 21088 17119 21140 17128
rect 21088 17085 21097 17119
rect 21097 17085 21131 17119
rect 21131 17085 21140 17119
rect 21088 17076 21140 17085
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 23020 17119 23072 17128
rect 23020 17085 23029 17119
rect 23029 17085 23063 17119
rect 23063 17085 23072 17119
rect 23020 17076 23072 17085
rect 20536 17008 20588 17060
rect 22192 17008 22244 17060
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 24032 17187 24084 17196
rect 24032 17153 24066 17187
rect 24066 17153 24084 17187
rect 24032 17144 24084 17153
rect 24768 17076 24820 17128
rect 25780 17051 25832 17060
rect 25780 17017 25789 17051
rect 25789 17017 25823 17051
rect 25823 17017 25832 17051
rect 25780 17008 25832 17017
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 14556 16940 14608 16992
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 20812 16983 20864 16992
rect 20812 16949 20821 16983
rect 20821 16949 20855 16983
rect 20855 16949 20864 16983
rect 20812 16940 20864 16949
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21824 16940 21876 16992
rect 22468 16940 22520 16992
rect 23296 16940 23348 16992
rect 23572 16940 23624 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 15936 16736 15988 16788
rect 18512 16736 18564 16788
rect 20260 16736 20312 16788
rect 5632 16668 5684 16720
rect 6644 16711 6696 16720
rect 6644 16677 6653 16711
rect 6653 16677 6687 16711
rect 6687 16677 6696 16711
rect 6644 16668 6696 16677
rect 22100 16668 22152 16720
rect 12256 16643 12308 16652
rect 12256 16609 12265 16643
rect 12265 16609 12299 16643
rect 12299 16609 12308 16643
rect 12256 16600 12308 16609
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 12440 16600 12492 16652
rect 13636 16600 13688 16652
rect 15200 16600 15252 16652
rect 15292 16600 15344 16652
rect 16856 16600 16908 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 18328 16600 18380 16652
rect 20904 16600 20956 16652
rect 18696 16532 18748 16584
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 1584 16396 1636 16448
rect 11612 16396 11664 16448
rect 12992 16464 13044 16516
rect 19156 16464 19208 16516
rect 19708 16464 19760 16516
rect 20904 16464 20956 16516
rect 21272 16464 21324 16516
rect 21824 16575 21876 16584
rect 21824 16541 21833 16575
rect 21833 16541 21867 16575
rect 21867 16541 21876 16575
rect 21824 16532 21876 16541
rect 21916 16507 21968 16516
rect 21916 16473 21925 16507
rect 21925 16473 21959 16507
rect 21959 16473 21968 16507
rect 21916 16464 21968 16473
rect 23020 16532 23072 16584
rect 12808 16396 12860 16448
rect 12900 16439 12952 16448
rect 12900 16405 12909 16439
rect 12909 16405 12943 16439
rect 12943 16405 12952 16439
rect 12900 16396 12952 16405
rect 15844 16439 15896 16448
rect 15844 16405 15853 16439
rect 15853 16405 15887 16439
rect 15887 16405 15896 16439
rect 15844 16396 15896 16405
rect 21088 16396 21140 16448
rect 21548 16439 21600 16448
rect 21548 16405 21557 16439
rect 21557 16405 21591 16439
rect 21591 16405 21600 16439
rect 21548 16396 21600 16405
rect 21732 16396 21784 16448
rect 23756 16439 23808 16448
rect 23756 16405 23765 16439
rect 23765 16405 23799 16439
rect 23799 16405 23808 16439
rect 23756 16396 23808 16405
rect 23848 16439 23900 16448
rect 23848 16405 23857 16439
rect 23857 16405 23891 16439
rect 23891 16405 23900 16439
rect 23848 16396 23900 16405
rect 25504 16396 25556 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 4620 16192 4672 16244
rect 5816 16192 5868 16244
rect 12440 16192 12492 16244
rect 18328 16235 18380 16244
rect 18328 16201 18337 16235
rect 18337 16201 18371 16235
rect 18371 16201 18380 16235
rect 18328 16192 18380 16201
rect 1768 16124 1820 16176
rect 848 16056 900 16108
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2412 16056 2464 16108
rect 3884 16056 3936 16108
rect 4804 16056 4856 16108
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 4712 15852 4764 15904
rect 5540 16124 5592 16176
rect 6184 16124 6236 16176
rect 11704 16124 11756 16176
rect 6368 16099 6420 16108
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 12072 16056 12124 16108
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 20812 16192 20864 16244
rect 23756 16192 23808 16244
rect 23848 16192 23900 16244
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 19708 16099 19760 16108
rect 19708 16065 19726 16099
rect 19726 16065 19760 16099
rect 19708 16056 19760 16065
rect 10968 15988 11020 16040
rect 13636 16031 13688 16040
rect 13636 15997 13645 16031
rect 13645 15997 13679 16031
rect 13679 15997 13688 16031
rect 13636 15988 13688 15997
rect 5908 15963 5960 15972
rect 5908 15929 5917 15963
rect 5917 15929 5951 15963
rect 5951 15929 5960 15963
rect 5908 15920 5960 15929
rect 6552 15852 6604 15904
rect 11796 15852 11848 15904
rect 12256 15852 12308 15904
rect 20904 16056 20956 16108
rect 21548 16056 21600 16108
rect 23020 16124 23072 16176
rect 21732 15988 21784 16040
rect 15292 15852 15344 15904
rect 17868 15852 17920 15904
rect 18696 15852 18748 15904
rect 20260 15895 20312 15904
rect 20260 15861 20269 15895
rect 20269 15861 20303 15895
rect 20303 15861 20312 15895
rect 20260 15852 20312 15861
rect 20352 15852 20404 15904
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 22100 16056 22152 16108
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 22652 16099 22704 16108
rect 22652 16065 22661 16099
rect 22661 16065 22695 16099
rect 22695 16065 22704 16099
rect 22652 16056 22704 16065
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 23572 16099 23624 16108
rect 23572 16065 23581 16099
rect 23581 16065 23615 16099
rect 23615 16065 23624 16099
rect 23572 16056 23624 16065
rect 23848 16099 23900 16108
rect 23848 16065 23857 16099
rect 23857 16065 23891 16099
rect 23891 16065 23900 16099
rect 23848 16056 23900 16065
rect 25504 16099 25556 16108
rect 25504 16065 25513 16099
rect 25513 16065 25547 16099
rect 25547 16065 25556 16099
rect 25504 16056 25556 16065
rect 25688 16056 25740 16108
rect 22652 15920 22704 15972
rect 23112 15920 23164 15972
rect 24492 15920 24544 15972
rect 24768 15963 24820 15972
rect 24768 15929 24777 15963
rect 24777 15929 24811 15963
rect 24811 15929 24820 15963
rect 24768 15920 24820 15929
rect 24584 15852 24636 15904
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 1768 15648 1820 15700
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 2596 15691 2648 15700
rect 2596 15657 2605 15691
rect 2605 15657 2639 15691
rect 2639 15657 2648 15691
rect 2596 15648 2648 15657
rect 6736 15648 6788 15700
rect 11704 15648 11756 15700
rect 12072 15648 12124 15700
rect 13360 15648 13412 15700
rect 21364 15648 21416 15700
rect 23756 15648 23808 15700
rect 26056 15648 26108 15700
rect 12808 15580 12860 15632
rect 3240 15512 3292 15564
rect 3332 15512 3384 15564
rect 1492 15419 1544 15428
rect 1492 15385 1501 15419
rect 1501 15385 1535 15419
rect 1535 15385 1544 15419
rect 1492 15376 1544 15385
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 3608 15444 3660 15496
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 2688 15376 2740 15428
rect 3332 15419 3384 15428
rect 3332 15385 3341 15419
rect 3341 15385 3375 15419
rect 3375 15385 3384 15419
rect 3332 15376 3384 15385
rect 3976 15419 4028 15428
rect 3976 15385 3985 15419
rect 3985 15385 4019 15419
rect 4019 15385 4028 15419
rect 3976 15376 4028 15385
rect 5908 15512 5960 15564
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 7380 15444 7432 15496
rect 8576 15444 8628 15496
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 13636 15512 13688 15564
rect 9036 15376 9088 15428
rect 9588 15376 9640 15428
rect 12256 15444 12308 15496
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 13176 15444 13228 15496
rect 15292 15512 15344 15564
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 18512 15580 18564 15632
rect 20352 15580 20404 15632
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 22652 15580 22704 15632
rect 17960 15512 18012 15521
rect 21732 15512 21784 15564
rect 22744 15512 22796 15564
rect 24952 15555 25004 15564
rect 24952 15521 24961 15555
rect 24961 15521 24995 15555
rect 24995 15521 25004 15555
rect 24952 15512 25004 15521
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 3148 15351 3200 15360
rect 3148 15317 3157 15351
rect 3157 15317 3191 15351
rect 3191 15317 3200 15351
rect 3148 15308 3200 15317
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 4804 15308 4856 15360
rect 5356 15351 5408 15360
rect 5356 15317 5365 15351
rect 5365 15317 5399 15351
rect 5399 15317 5408 15351
rect 5356 15308 5408 15317
rect 6736 15308 6788 15360
rect 8944 15308 8996 15360
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 13636 15419 13688 15428
rect 13636 15385 13645 15419
rect 13645 15385 13679 15419
rect 13679 15385 13688 15419
rect 13636 15376 13688 15385
rect 18512 15376 18564 15428
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 20168 15444 20220 15496
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 21916 15487 21968 15496
rect 21916 15453 21925 15487
rect 21925 15453 21959 15487
rect 21959 15453 21968 15487
rect 21916 15444 21968 15453
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 23664 15444 23716 15496
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 20260 15376 20312 15428
rect 23296 15376 23348 15428
rect 23388 15376 23440 15428
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 15936 15351 15988 15360
rect 15936 15317 15945 15351
rect 15945 15317 15979 15351
rect 15979 15317 15988 15351
rect 15936 15308 15988 15317
rect 18604 15351 18656 15360
rect 18604 15317 18613 15351
rect 18613 15317 18647 15351
rect 18647 15317 18656 15351
rect 18604 15308 18656 15317
rect 20996 15308 21048 15360
rect 24308 15308 24360 15360
rect 25412 15351 25464 15360
rect 25412 15317 25421 15351
rect 25421 15317 25455 15351
rect 25455 15317 25464 15351
rect 25412 15308 25464 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 3148 15104 3200 15156
rect 3976 15104 4028 15156
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 2872 14968 2924 15020
rect 3148 14968 3200 15020
rect 4160 14968 4212 15020
rect 1860 14764 1912 14816
rect 3056 14943 3108 14952
rect 3056 14909 3065 14943
rect 3065 14909 3099 14943
rect 3099 14909 3108 14943
rect 3056 14900 3108 14909
rect 5540 15104 5592 15156
rect 13268 15104 13320 15156
rect 13360 15104 13412 15156
rect 5356 15036 5408 15088
rect 5816 15036 5868 15088
rect 6000 14968 6052 15020
rect 6644 14968 6696 15020
rect 7656 14968 7708 15020
rect 5724 14900 5776 14952
rect 2688 14832 2740 14884
rect 6644 14875 6696 14884
rect 6644 14841 6653 14875
rect 6653 14841 6687 14875
rect 6687 14841 6696 14875
rect 6644 14832 6696 14841
rect 9128 14968 9180 15020
rect 9220 14968 9272 15020
rect 9772 14968 9824 15020
rect 10968 15036 11020 15088
rect 12348 15036 12400 15088
rect 10232 15011 10284 15020
rect 10232 14977 10266 15011
rect 10266 14977 10284 15011
rect 10232 14968 10284 14977
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 13084 14968 13136 15020
rect 13360 15011 13412 15020
rect 13360 14977 13378 15011
rect 13378 14977 13412 15011
rect 13360 14968 13412 14977
rect 14004 15011 14056 15020
rect 14004 14977 14038 15011
rect 14038 14977 14056 15011
rect 14004 14968 14056 14977
rect 15200 14900 15252 14952
rect 15936 15104 15988 15156
rect 22008 15104 22060 15156
rect 15752 15036 15804 15088
rect 17132 15036 17184 15088
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 21456 14968 21508 15020
rect 23296 15147 23348 15156
rect 23296 15113 23305 15147
rect 23305 15113 23339 15147
rect 23339 15113 23348 15147
rect 23296 15104 23348 15113
rect 24308 15104 24360 15156
rect 25228 15104 25280 15156
rect 23756 15079 23808 15088
rect 23756 15045 23765 15079
rect 23765 15045 23799 15079
rect 23799 15045 23808 15079
rect 23756 15036 23808 15045
rect 24952 15011 25004 15020
rect 24952 14977 24961 15011
rect 24961 14977 24995 15011
rect 24995 14977 25004 15011
rect 24952 14968 25004 14977
rect 15568 14832 15620 14884
rect 16764 14900 16816 14952
rect 20444 14900 20496 14952
rect 17316 14832 17368 14884
rect 22652 14832 22704 14884
rect 2872 14764 2924 14816
rect 3332 14764 3384 14816
rect 3700 14764 3752 14816
rect 4988 14764 5040 14816
rect 5632 14764 5684 14816
rect 6092 14764 6144 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 13912 14764 13964 14816
rect 14832 14764 14884 14816
rect 15384 14764 15436 14816
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 21732 14764 21784 14816
rect 24860 14764 24912 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 3240 14603 3292 14612
rect 3240 14569 3249 14603
rect 3249 14569 3283 14603
rect 3283 14569 3292 14603
rect 3240 14560 3292 14569
rect 3424 14560 3476 14612
rect 3700 14560 3752 14612
rect 3332 14492 3384 14544
rect 4804 14560 4856 14612
rect 5080 14560 5132 14612
rect 3148 14424 3200 14476
rect 1584 14356 1636 14408
rect 3056 14356 3108 14408
rect 8116 14560 8168 14612
rect 9588 14560 9640 14612
rect 11612 14560 11664 14612
rect 17316 14560 17368 14612
rect 18604 14560 18656 14612
rect 5264 14492 5316 14544
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 3700 14356 3752 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 2136 14288 2188 14340
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 4804 14356 4856 14408
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 5356 14424 5408 14476
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 5540 14356 5592 14408
rect 6184 14356 6236 14408
rect 6552 14356 6604 14408
rect 6644 14356 6696 14408
rect 8024 14356 8076 14408
rect 8576 14356 8628 14408
rect 11980 14492 12032 14544
rect 17132 14535 17184 14544
rect 17132 14501 17141 14535
rect 17141 14501 17175 14535
rect 17175 14501 17184 14535
rect 17132 14492 17184 14501
rect 11336 14424 11388 14476
rect 12164 14424 12216 14476
rect 5816 14288 5868 14340
rect 9772 14356 9824 14408
rect 11796 14356 11848 14408
rect 11980 14356 12032 14408
rect 12992 14467 13044 14476
rect 12992 14433 13001 14467
rect 13001 14433 13035 14467
rect 13035 14433 13044 14467
rect 12992 14424 13044 14433
rect 13912 14467 13964 14476
rect 13912 14433 13921 14467
rect 13921 14433 13955 14467
rect 13955 14433 13964 14467
rect 13912 14424 13964 14433
rect 20260 14560 20312 14612
rect 22192 14560 22244 14612
rect 22836 14560 22888 14612
rect 20812 14492 20864 14544
rect 12624 14288 12676 14340
rect 15200 14288 15252 14340
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16948 14356 17000 14408
rect 18512 14356 18564 14408
rect 16672 14288 16724 14340
rect 18604 14288 18656 14340
rect 20444 14288 20496 14340
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 6460 14220 6512 14272
rect 7472 14220 7524 14272
rect 9312 14220 9364 14272
rect 9588 14220 9640 14272
rect 12348 14220 12400 14272
rect 13544 14220 13596 14272
rect 15292 14220 15344 14272
rect 15384 14220 15436 14272
rect 18972 14220 19024 14272
rect 19800 14220 19852 14272
rect 20720 14220 20772 14272
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 23388 14356 23440 14408
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 21824 14331 21876 14340
rect 21824 14297 21833 14331
rect 21833 14297 21867 14331
rect 21867 14297 21876 14331
rect 21824 14288 21876 14297
rect 24308 14288 24360 14340
rect 23204 14220 23256 14272
rect 24032 14220 24084 14272
rect 25688 14220 25740 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 112 14016 164 14068
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 1860 13923 1912 13932
rect 1860 13889 1894 13923
rect 1894 13889 1912 13923
rect 1860 13880 1912 13889
rect 2964 13880 3016 13932
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 5264 13948 5316 14000
rect 2872 13812 2924 13864
rect 3148 13812 3200 13864
rect 3792 13880 3844 13932
rect 4804 13880 4856 13932
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 4988 13719 5040 13728
rect 4988 13685 4997 13719
rect 4997 13685 5031 13719
rect 5031 13685 5040 13719
rect 4988 13676 5040 13685
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 6276 13948 6328 14000
rect 6460 13948 6512 14000
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6000 13880 6052 13932
rect 8024 13991 8076 14000
rect 8024 13957 8033 13991
rect 8033 13957 8067 13991
rect 8067 13957 8076 13991
rect 8024 13948 8076 13957
rect 8300 13948 8352 14000
rect 5356 13744 5408 13796
rect 5632 13744 5684 13796
rect 6000 13744 6052 13796
rect 6644 13812 6696 13864
rect 7472 13880 7524 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 8760 13948 8812 14000
rect 9404 13991 9456 14000
rect 9404 13957 9413 13991
rect 9413 13957 9447 13991
rect 9447 13957 9456 13991
rect 9404 13948 9456 13957
rect 9496 13948 9548 14000
rect 7748 13880 7800 13889
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 8116 13744 8168 13796
rect 8484 13812 8536 13864
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 5816 13676 5868 13728
rect 7840 13676 7892 13728
rect 8300 13676 8352 13728
rect 9128 13880 9180 13932
rect 9312 13880 9364 13932
rect 12164 13991 12216 14000
rect 12164 13957 12173 13991
rect 12173 13957 12207 13991
rect 12207 13957 12216 13991
rect 12164 13948 12216 13957
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 15844 14016 15896 14068
rect 16212 14016 16264 14068
rect 18512 14059 18564 14068
rect 18512 14025 18521 14059
rect 18521 14025 18555 14059
rect 18555 14025 18564 14059
rect 18512 14016 18564 14025
rect 18604 14059 18656 14068
rect 18604 14025 18613 14059
rect 18613 14025 18647 14059
rect 18647 14025 18656 14059
rect 18604 14016 18656 14025
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 15384 13991 15436 14000
rect 15384 13957 15396 13991
rect 15396 13957 15436 13991
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 11796 13923 11848 13932
rect 11796 13889 11805 13923
rect 11805 13889 11839 13923
rect 11839 13889 11848 13923
rect 11796 13880 11848 13889
rect 15384 13948 15436 13957
rect 19800 14059 19852 14068
rect 19800 14025 19809 14059
rect 19809 14025 19843 14059
rect 19843 14025 19852 14059
rect 19800 14016 19852 14025
rect 20076 14016 20128 14068
rect 21088 14016 21140 14068
rect 21364 14016 21416 14068
rect 23388 14016 23440 14068
rect 24308 14059 24360 14068
rect 24308 14025 24317 14059
rect 24317 14025 24351 14059
rect 24351 14025 24360 14059
rect 24308 14016 24360 14025
rect 25412 14059 25464 14068
rect 25412 14025 25421 14059
rect 25421 14025 25455 14059
rect 25455 14025 25464 14059
rect 25412 14016 25464 14025
rect 25780 14059 25832 14068
rect 25780 14025 25789 14059
rect 25789 14025 25823 14059
rect 25823 14025 25832 14059
rect 25780 14016 25832 14025
rect 12808 13880 12860 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 12624 13812 12676 13864
rect 13636 13812 13688 13864
rect 16856 13880 16908 13932
rect 16948 13880 17000 13932
rect 19524 13880 19576 13932
rect 20168 13880 20220 13932
rect 23756 13948 23808 14000
rect 20352 13880 20404 13932
rect 20904 13880 20956 13932
rect 21640 13880 21692 13932
rect 21916 13880 21968 13932
rect 24492 13948 24544 14000
rect 25688 13948 25740 14000
rect 18328 13744 18380 13796
rect 9036 13676 9088 13728
rect 9220 13676 9272 13728
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 11888 13676 11940 13728
rect 12072 13676 12124 13728
rect 12440 13676 12492 13728
rect 20444 13676 20496 13728
rect 21456 13744 21508 13796
rect 21732 13744 21784 13796
rect 24032 13923 24084 13932
rect 24032 13889 24041 13923
rect 24041 13889 24075 13923
rect 24075 13889 24084 13923
rect 24032 13880 24084 13889
rect 24124 13880 24176 13932
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 21548 13676 21600 13728
rect 22928 13676 22980 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2136 13515 2188 13524
rect 2136 13481 2145 13515
rect 2145 13481 2179 13515
rect 2179 13481 2188 13515
rect 2136 13472 2188 13481
rect 2596 13472 2648 13524
rect 5264 13472 5316 13524
rect 6276 13515 6328 13524
rect 6276 13481 6285 13515
rect 6285 13481 6319 13515
rect 6319 13481 6328 13515
rect 6276 13472 6328 13481
rect 7012 13472 7064 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 8024 13472 8076 13524
rect 8760 13472 8812 13524
rect 10048 13472 10100 13524
rect 14004 13472 14056 13524
rect 15384 13472 15436 13524
rect 18236 13472 18288 13524
rect 5448 13447 5500 13456
rect 5448 13413 5457 13447
rect 5457 13413 5491 13447
rect 5491 13413 5500 13447
rect 5448 13404 5500 13413
rect 6184 13404 6236 13456
rect 4988 13268 5040 13320
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 5724 13268 5776 13320
rect 8300 13336 8352 13388
rect 6828 13268 6880 13320
rect 2688 13200 2740 13252
rect 3332 13132 3384 13184
rect 7472 13268 7524 13320
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 9128 13336 9180 13388
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 8208 13200 8260 13252
rect 9496 13268 9548 13320
rect 8668 13200 8720 13252
rect 9588 13200 9640 13252
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 16212 13379 16264 13388
rect 16212 13345 16221 13379
rect 16221 13345 16255 13379
rect 16255 13345 16264 13379
rect 16212 13336 16264 13345
rect 16948 13336 17000 13388
rect 20352 13472 20404 13524
rect 20812 13472 20864 13524
rect 21088 13472 21140 13524
rect 21548 13472 21600 13524
rect 21916 13472 21968 13524
rect 19892 13404 19944 13456
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 18236 13268 18288 13320
rect 20260 13268 20312 13320
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 12992 13200 13044 13252
rect 14280 13200 14332 13252
rect 15292 13200 15344 13252
rect 17868 13200 17920 13252
rect 8024 13132 8076 13184
rect 8484 13132 8536 13184
rect 9312 13132 9364 13184
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 21548 13268 21600 13320
rect 23204 13404 23256 13456
rect 24124 13404 24176 13456
rect 23388 13268 23440 13320
rect 21180 13243 21232 13252
rect 21180 13209 21214 13243
rect 21214 13209 21232 13243
rect 21180 13200 21232 13209
rect 21824 13200 21876 13252
rect 21272 13132 21324 13184
rect 22100 13132 22152 13184
rect 22928 13200 22980 13252
rect 23204 13200 23256 13252
rect 22744 13175 22796 13184
rect 22744 13141 22753 13175
rect 22753 13141 22787 13175
rect 22787 13141 22796 13175
rect 22744 13132 22796 13141
rect 23664 13200 23716 13252
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 24032 13268 24084 13320
rect 24400 13311 24452 13320
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 24124 13200 24176 13252
rect 23940 13132 23992 13184
rect 25596 13132 25648 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 6184 12928 6236 12980
rect 7840 12928 7892 12980
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 5816 12860 5868 12912
rect 7748 12860 7800 12912
rect 8392 12928 8444 12980
rect 8668 12928 8720 12980
rect 8576 12860 8628 12912
rect 8944 12903 8996 12912
rect 8944 12869 8969 12903
rect 8969 12869 8996 12903
rect 17868 12971 17920 12980
rect 17868 12937 17877 12971
rect 17877 12937 17911 12971
rect 17911 12937 17920 12971
rect 17868 12928 17920 12937
rect 19248 12928 19300 12980
rect 19524 12971 19576 12980
rect 19524 12937 19533 12971
rect 19533 12937 19567 12971
rect 19567 12937 19576 12971
rect 19524 12928 19576 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 8944 12860 8996 12869
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 4620 12792 4672 12844
rect 4804 12724 4856 12776
rect 5448 12835 5500 12844
rect 5448 12801 5457 12835
rect 5457 12801 5491 12835
rect 5491 12801 5500 12835
rect 5448 12792 5500 12801
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 8024 12792 8076 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 12900 12792 12952 12844
rect 19616 12792 19668 12844
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 19892 12792 19944 12844
rect 6828 12724 6880 12776
rect 10968 12724 11020 12776
rect 18236 12724 18288 12776
rect 19064 12724 19116 12776
rect 19524 12724 19576 12776
rect 20444 12792 20496 12844
rect 5540 12656 5592 12708
rect 22744 12860 22796 12912
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 21180 12792 21232 12844
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 21640 12835 21692 12844
rect 21640 12801 21649 12835
rect 21649 12801 21683 12835
rect 21683 12801 21692 12835
rect 21640 12792 21692 12801
rect 24124 12928 24176 12980
rect 25780 12971 25832 12980
rect 25780 12937 25789 12971
rect 25789 12937 25823 12971
rect 25823 12937 25832 12971
rect 25780 12928 25832 12937
rect 23480 12860 23532 12912
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 23664 12835 23716 12844
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 23940 12835 23992 12844
rect 23940 12801 23949 12835
rect 23949 12801 23983 12835
rect 23983 12801 23992 12835
rect 23940 12792 23992 12801
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 25044 12792 25096 12844
rect 25596 12835 25648 12844
rect 25596 12801 25611 12835
rect 25611 12801 25645 12835
rect 25645 12801 25648 12835
rect 25596 12792 25648 12801
rect 22008 12724 22060 12776
rect 23756 12724 23808 12776
rect 3424 12588 3476 12640
rect 4712 12588 4764 12640
rect 7288 12588 7340 12640
rect 9312 12588 9364 12640
rect 13268 12588 13320 12640
rect 20720 12588 20772 12640
rect 25136 12588 25188 12640
rect 25412 12631 25464 12640
rect 25412 12597 25421 12631
rect 25421 12597 25455 12631
rect 25455 12597 25464 12631
rect 25412 12588 25464 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2596 12384 2648 12436
rect 3608 12316 3660 12368
rect 5632 12384 5684 12436
rect 8944 12427 8996 12436
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 19616 12384 19668 12436
rect 20168 12384 20220 12436
rect 2872 12248 2924 12300
rect 5632 12248 5684 12300
rect 7196 12248 7248 12300
rect 9036 12248 9088 12300
rect 1400 12112 1452 12164
rect 1952 12044 2004 12096
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 2688 12155 2740 12164
rect 2688 12121 2697 12155
rect 2697 12121 2731 12155
rect 2731 12121 2740 12155
rect 2688 12112 2740 12121
rect 2964 12155 3016 12164
rect 2964 12121 2973 12155
rect 2973 12121 3007 12155
rect 3007 12121 3016 12155
rect 2964 12112 3016 12121
rect 3148 12155 3200 12164
rect 3148 12121 3157 12155
rect 3157 12121 3191 12155
rect 3191 12121 3200 12155
rect 3424 12155 3476 12164
rect 3148 12112 3200 12121
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 3424 12121 3446 12155
rect 3446 12121 3476 12155
rect 3424 12112 3476 12121
rect 4436 12180 4488 12232
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 8300 12223 8352 12232
rect 8300 12189 8309 12223
rect 8309 12189 8343 12223
rect 8343 12189 8352 12223
rect 8300 12180 8352 12189
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 5264 12112 5316 12164
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 9496 12248 9548 12300
rect 10968 12248 11020 12300
rect 8760 12180 8812 12189
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 13084 12248 13136 12300
rect 3700 12044 3752 12096
rect 3792 12044 3844 12096
rect 4068 12044 4120 12096
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 5816 12044 5868 12096
rect 6736 12044 6788 12096
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 13360 12180 13412 12232
rect 14740 12180 14792 12232
rect 14832 12180 14884 12232
rect 16856 12248 16908 12300
rect 19800 12248 19852 12300
rect 14556 12112 14608 12164
rect 14188 12044 14240 12096
rect 14464 12044 14516 12096
rect 15568 12044 15620 12096
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 16580 12044 16632 12096
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 19708 12180 19760 12232
rect 20260 12248 20312 12300
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20720 12316 20772 12368
rect 20536 12180 20588 12232
rect 21456 12316 21508 12368
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21824 12180 21876 12232
rect 23572 12384 23624 12436
rect 24768 12384 24820 12436
rect 25044 12427 25096 12436
rect 25044 12393 25053 12427
rect 25053 12393 25087 12427
rect 25087 12393 25096 12427
rect 25044 12384 25096 12393
rect 25136 12427 25188 12436
rect 25136 12393 25145 12427
rect 25145 12393 25179 12427
rect 25179 12393 25188 12427
rect 25136 12384 25188 12393
rect 23480 12316 23532 12368
rect 24400 12316 24452 12368
rect 23848 12248 23900 12300
rect 24308 12248 24360 12300
rect 24492 12248 24544 12300
rect 22652 12180 22704 12232
rect 23388 12180 23440 12232
rect 19340 12044 19392 12096
rect 20168 12044 20220 12096
rect 20444 12044 20496 12096
rect 22100 12044 22152 12096
rect 22928 12112 22980 12164
rect 24676 12223 24728 12232
rect 24676 12189 24685 12223
rect 24685 12189 24719 12223
rect 24719 12189 24728 12223
rect 24676 12180 24728 12189
rect 24860 12180 24912 12232
rect 25688 12223 25740 12232
rect 25688 12189 25697 12223
rect 25697 12189 25731 12223
rect 25731 12189 25740 12223
rect 25688 12180 25740 12189
rect 23204 12044 23256 12096
rect 25412 12155 25464 12164
rect 25412 12121 25421 12155
rect 25421 12121 25455 12155
rect 25455 12121 25464 12155
rect 25412 12112 25464 12121
rect 25596 12044 25648 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2412 11840 2464 11892
rect 2872 11840 2924 11892
rect 3700 11840 3752 11892
rect 3976 11840 4028 11892
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 3056 11772 3108 11824
rect 3424 11772 3476 11824
rect 1952 11747 2004 11756
rect 1952 11713 1986 11747
rect 1986 11713 2004 11747
rect 1952 11704 2004 11713
rect 3884 11815 3936 11824
rect 3884 11781 3893 11815
rect 3893 11781 3927 11815
rect 3927 11781 3936 11815
rect 4804 11840 4856 11892
rect 5264 11840 5316 11892
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 8484 11840 8536 11892
rect 12440 11840 12492 11892
rect 3884 11772 3936 11781
rect 4436 11772 4488 11824
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 8760 11772 8812 11824
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 14556 11840 14608 11892
rect 19340 11840 19392 11892
rect 21364 11840 21416 11892
rect 25780 11883 25832 11892
rect 25780 11849 25789 11883
rect 25789 11849 25823 11883
rect 25823 11849 25832 11883
rect 25780 11840 25832 11849
rect 4804 11636 4856 11688
rect 3608 11611 3660 11620
rect 3608 11577 3617 11611
rect 3617 11577 3651 11611
rect 3651 11577 3660 11611
rect 3608 11568 3660 11577
rect 4712 11568 4764 11620
rect 5172 11747 5224 11756
rect 5172 11713 5181 11747
rect 5181 11713 5215 11747
rect 5215 11713 5224 11747
rect 5172 11704 5224 11713
rect 5264 11704 5316 11756
rect 5356 11636 5408 11688
rect 6736 11704 6788 11756
rect 7840 11704 7892 11756
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 8852 11704 8904 11756
rect 10968 11704 11020 11756
rect 11796 11747 11848 11756
rect 11796 11713 11830 11747
rect 11830 11713 11848 11747
rect 11796 11704 11848 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 8208 11636 8260 11688
rect 13176 11568 13228 11620
rect 2964 11500 3016 11552
rect 3884 11500 3936 11552
rect 4620 11500 4672 11552
rect 4804 11500 4856 11552
rect 5632 11500 5684 11552
rect 8944 11500 8996 11552
rect 13636 11815 13688 11824
rect 13636 11781 13645 11815
rect 13645 11781 13679 11815
rect 13679 11781 13688 11815
rect 13636 11772 13688 11781
rect 17316 11815 17368 11824
rect 17316 11781 17350 11815
rect 17350 11781 17368 11815
rect 17316 11772 17368 11781
rect 13912 11704 13964 11756
rect 14464 11704 14516 11756
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 15568 11704 15620 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 19248 11704 19300 11756
rect 20904 11772 20956 11824
rect 19892 11747 19944 11756
rect 19892 11713 19926 11747
rect 19926 11713 19944 11747
rect 19892 11704 19944 11713
rect 20168 11704 20220 11756
rect 23664 11772 23716 11824
rect 24584 11772 24636 11824
rect 21916 11704 21968 11756
rect 24124 11747 24176 11756
rect 24124 11713 24158 11747
rect 24158 11713 24176 11747
rect 24124 11704 24176 11713
rect 14188 11679 14240 11688
rect 14188 11645 14197 11679
rect 14197 11645 14231 11679
rect 14231 11645 14240 11679
rect 14188 11636 14240 11645
rect 14188 11500 14240 11552
rect 18972 11679 19024 11688
rect 18972 11645 18981 11679
rect 18981 11645 19015 11679
rect 19015 11645 19024 11679
rect 18972 11636 19024 11645
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 20720 11568 20772 11620
rect 21824 11568 21876 11620
rect 15660 11500 15712 11552
rect 16028 11500 16080 11552
rect 16580 11500 16632 11552
rect 17408 11500 17460 11552
rect 18512 11543 18564 11552
rect 18512 11509 18521 11543
rect 18521 11509 18555 11543
rect 18555 11509 18564 11543
rect 18512 11500 18564 11509
rect 20536 11500 20588 11552
rect 22100 11500 22152 11552
rect 23664 11568 23716 11620
rect 25596 11747 25648 11756
rect 25596 11713 25605 11747
rect 25605 11713 25639 11747
rect 25639 11713 25648 11747
rect 25596 11704 25648 11713
rect 25596 11568 25648 11620
rect 23204 11543 23256 11552
rect 23204 11509 23213 11543
rect 23213 11509 23247 11543
rect 23247 11509 23256 11543
rect 23204 11500 23256 11509
rect 25320 11500 25372 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4804 11296 4856 11348
rect 5540 11296 5592 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 3056 11092 3108 11144
rect 3240 11024 3292 11076
rect 3792 11067 3844 11076
rect 3792 11033 3801 11067
rect 3801 11033 3835 11067
rect 3835 11033 3844 11067
rect 3792 11024 3844 11033
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4712 11160 4764 11212
rect 5264 11092 5316 11144
rect 7288 11296 7340 11348
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 8300 11296 8352 11348
rect 8484 11228 8536 11280
rect 8852 11296 8904 11348
rect 11796 11296 11848 11348
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 14188 11296 14240 11348
rect 8944 11228 8996 11280
rect 8024 11160 8076 11212
rect 4344 11024 4396 11076
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 5724 11024 5776 11076
rect 6736 11024 6788 11076
rect 4160 10999 4212 11008
rect 4160 10965 4169 10999
rect 4169 10965 4203 10999
rect 4203 10965 4212 10999
rect 4160 10956 4212 10965
rect 7196 11067 7248 11076
rect 7196 11033 7205 11067
rect 7205 11033 7239 11067
rect 7239 11033 7248 11067
rect 7196 11024 7248 11033
rect 7380 11067 7432 11076
rect 7380 11033 7405 11067
rect 7405 11033 7432 11067
rect 7380 11024 7432 11033
rect 7656 11067 7708 11076
rect 7656 11033 7665 11067
rect 7665 11033 7699 11067
rect 7699 11033 7708 11067
rect 7656 11024 7708 11033
rect 8576 11160 8628 11212
rect 13084 11228 13136 11280
rect 14832 11296 14884 11348
rect 14924 11228 14976 11280
rect 18420 11296 18472 11348
rect 13268 11160 13320 11212
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 8668 11024 8720 11076
rect 12072 11024 12124 11076
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 8024 10956 8076 11008
rect 13636 11092 13688 11144
rect 14740 11160 14792 11212
rect 17040 11160 17092 11212
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19892 11296 19944 11348
rect 21916 11296 21968 11348
rect 22928 11296 22980 11348
rect 18972 11228 19024 11280
rect 20536 11160 20588 11212
rect 18512 11092 18564 11144
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 14556 11024 14608 11076
rect 15384 11024 15436 11076
rect 17408 11024 17460 11076
rect 20444 11135 20496 11144
rect 20444 11101 20453 11135
rect 20453 11101 20487 11135
rect 20487 11101 20496 11135
rect 20444 11092 20496 11101
rect 21364 11160 21416 11212
rect 22192 11228 22244 11280
rect 23572 11228 23624 11280
rect 21180 11135 21232 11144
rect 21180 11101 21189 11135
rect 21189 11101 21223 11135
rect 21223 11101 21232 11135
rect 21180 11092 21232 11101
rect 21456 11092 21508 11144
rect 21548 11092 21600 11144
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 23204 11160 23256 11212
rect 23388 11160 23440 11212
rect 23664 11160 23716 11212
rect 25780 11339 25832 11348
rect 25780 11305 25789 11339
rect 25789 11305 25823 11339
rect 25823 11305 25832 11339
rect 25780 11296 25832 11305
rect 14924 10956 14976 11008
rect 15936 10956 15988 11008
rect 17132 10956 17184 11008
rect 21824 11024 21876 11076
rect 22928 11024 22980 11076
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 24124 11092 24176 11144
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 24584 11024 24636 11033
rect 24860 11024 24912 11076
rect 25320 11092 25372 11144
rect 20628 10956 20680 11008
rect 20996 10956 21048 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3608 10752 3660 10804
rect 3792 10752 3844 10804
rect 3056 10684 3108 10736
rect 4160 10616 4212 10668
rect 4344 10684 4396 10736
rect 5724 10752 5776 10804
rect 7472 10752 7524 10804
rect 5540 10684 5592 10736
rect 7104 10684 7156 10736
rect 7656 10752 7708 10804
rect 12348 10752 12400 10804
rect 13176 10752 13228 10804
rect 14924 10752 14976 10804
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 16488 10752 16540 10804
rect 20076 10752 20128 10804
rect 8484 10684 8536 10736
rect 10968 10727 11020 10736
rect 10968 10693 10977 10727
rect 10977 10693 11011 10727
rect 11011 10693 11020 10727
rect 10968 10684 11020 10693
rect 9680 10616 9732 10668
rect 14648 10684 14700 10736
rect 16672 10684 16724 10736
rect 21548 10752 21600 10804
rect 22284 10752 22336 10804
rect 22652 10752 22704 10804
rect 23664 10752 23716 10804
rect 24676 10752 24728 10804
rect 25780 10795 25832 10804
rect 25780 10761 25789 10795
rect 25789 10761 25823 10795
rect 25823 10761 25832 10795
rect 25780 10752 25832 10761
rect 11244 10616 11296 10668
rect 6736 10591 6788 10600
rect 6736 10557 6745 10591
rect 6745 10557 6779 10591
rect 6779 10557 6788 10591
rect 6736 10548 6788 10557
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 13728 10548 13780 10600
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 17132 10616 17184 10668
rect 18972 10616 19024 10668
rect 23296 10684 23348 10736
rect 12072 10480 12124 10532
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 15660 10548 15712 10600
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 19064 10548 19116 10600
rect 21916 10548 21968 10600
rect 22376 10616 22428 10668
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 23756 10659 23808 10668
rect 23756 10625 23765 10659
rect 23765 10625 23799 10659
rect 23799 10625 23808 10659
rect 23756 10616 23808 10625
rect 24216 10616 24268 10668
rect 19984 10480 20036 10532
rect 20260 10480 20312 10532
rect 23756 10480 23808 10532
rect 23848 10480 23900 10532
rect 16396 10412 16448 10464
rect 17868 10412 17920 10464
rect 20996 10455 21048 10464
rect 20996 10421 21005 10455
rect 21005 10421 21039 10455
rect 21039 10421 21048 10455
rect 20996 10412 21048 10421
rect 24860 10412 24912 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12256 10208 12308 10260
rect 14188 10251 14240 10260
rect 14188 10217 14197 10251
rect 14197 10217 14231 10251
rect 14231 10217 14240 10251
rect 14188 10208 14240 10217
rect 14556 10208 14608 10260
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 21548 10208 21600 10260
rect 25780 10251 25832 10260
rect 25780 10217 25789 10251
rect 25789 10217 25823 10251
rect 25823 10217 25832 10251
rect 25780 10208 25832 10217
rect 3056 10004 3108 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 11244 10072 11296 10124
rect 22284 10183 22336 10192
rect 22284 10149 22293 10183
rect 22293 10149 22327 10183
rect 22327 10149 22336 10183
rect 22284 10140 22336 10149
rect 4712 10004 4764 10013
rect 10968 10004 11020 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 13728 10004 13780 10056
rect 11060 9936 11112 9988
rect 12440 9936 12492 9988
rect 9680 9868 9732 9920
rect 9956 9868 10008 9920
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 14556 10004 14608 10056
rect 19800 10115 19852 10124
rect 19800 10081 19809 10115
rect 19809 10081 19843 10115
rect 19843 10081 19852 10115
rect 19800 10072 19852 10081
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 17592 10047 17644 10056
rect 17592 10013 17601 10047
rect 17601 10013 17635 10047
rect 17635 10013 17644 10047
rect 17592 10004 17644 10013
rect 17868 10047 17920 10056
rect 17868 10013 17902 10047
rect 17902 10013 17920 10047
rect 17868 10004 17920 10013
rect 18420 10004 18472 10056
rect 18788 10004 18840 10056
rect 15200 9936 15252 9988
rect 15660 9936 15712 9988
rect 17500 9936 17552 9988
rect 14648 9868 14700 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 16488 9868 16540 9920
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 20628 10047 20680 10056
rect 20628 10013 20637 10047
rect 20637 10013 20671 10047
rect 20671 10013 20680 10047
rect 20628 10004 20680 10013
rect 20996 10004 21048 10056
rect 24032 10004 24084 10056
rect 24768 10072 24820 10124
rect 24860 10004 24912 10056
rect 25136 10004 25188 10056
rect 22468 9936 22520 9988
rect 23940 9936 23992 9988
rect 24400 9936 24452 9988
rect 21272 9868 21324 9920
rect 23480 9868 23532 9920
rect 25596 10047 25648 10056
rect 25596 10013 25605 10047
rect 25605 10013 25639 10047
rect 25639 10013 25648 10047
rect 25596 10004 25648 10013
rect 25412 9911 25464 9920
rect 25412 9877 25421 9911
rect 25421 9877 25455 9911
rect 25455 9877 25464 9911
rect 25412 9868 25464 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1768 9596 1820 9648
rect 2596 9460 2648 9512
rect 12164 9596 12216 9648
rect 15108 9596 15160 9648
rect 15384 9596 15436 9648
rect 16396 9596 16448 9648
rect 10232 9571 10284 9580
rect 10232 9537 10266 9571
rect 10266 9537 10284 9571
rect 2964 9392 3016 9444
rect 10232 9528 10284 9537
rect 10968 9528 11020 9580
rect 14740 9528 14792 9580
rect 9588 9460 9640 9512
rect 4896 9392 4948 9444
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 16488 9460 16540 9512
rect 19248 9596 19300 9648
rect 22376 9664 22428 9716
rect 20076 9596 20128 9648
rect 18972 9528 19024 9580
rect 20168 9528 20220 9580
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 16580 9392 16632 9444
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 17592 9460 17644 9469
rect 2780 9324 2832 9376
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 3424 9324 3476 9376
rect 4804 9324 4856 9376
rect 6552 9324 6604 9376
rect 11060 9324 11112 9376
rect 12164 9324 12216 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13728 9324 13780 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 16488 9324 16540 9376
rect 20628 9460 20680 9512
rect 22008 9460 22060 9512
rect 23664 9528 23716 9580
rect 23848 9571 23900 9580
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 19340 9392 19392 9444
rect 17776 9324 17828 9376
rect 19984 9324 20036 9376
rect 20444 9324 20496 9376
rect 20812 9324 20864 9376
rect 25228 9367 25280 9376
rect 25228 9333 25237 9367
rect 25237 9333 25271 9367
rect 25271 9333 25280 9367
rect 25228 9324 25280 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1952 9120 2004 9172
rect 2780 8959 2832 8968
rect 2780 8925 2798 8959
rect 2798 8925 2832 8959
rect 2780 8916 2832 8925
rect 2964 8916 3016 8968
rect 3516 9120 3568 9172
rect 3608 9052 3660 9104
rect 4712 8916 4764 8968
rect 5448 9120 5500 9172
rect 6460 9120 6512 9172
rect 5908 9052 5960 9104
rect 6184 9052 6236 9104
rect 7196 9095 7248 9104
rect 7196 9061 7205 9095
rect 7205 9061 7239 9095
rect 7239 9061 7248 9095
rect 7196 9052 7248 9061
rect 7932 9052 7984 9104
rect 6552 8984 6604 9036
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 4620 8848 4672 8900
rect 4896 8891 4948 8900
rect 4896 8857 4905 8891
rect 4905 8857 4939 8891
rect 4939 8857 4948 8891
rect 4896 8848 4948 8857
rect 5540 8848 5592 8900
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 5908 8848 5960 8900
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 9956 9120 10008 9172
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 12900 9120 12952 9172
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 18972 9120 19024 9172
rect 11520 8916 11572 8968
rect 3424 8780 3476 8832
rect 4712 8780 4764 8832
rect 5724 8780 5776 8832
rect 6736 8780 6788 8832
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 10508 8848 10560 8900
rect 13636 8916 13688 8968
rect 13820 8916 13872 8968
rect 14740 8984 14792 9036
rect 17684 8984 17736 9036
rect 19616 8984 19668 9036
rect 20536 8984 20588 9036
rect 16488 8916 16540 8968
rect 19340 8916 19392 8968
rect 10232 8780 10284 8832
rect 11244 8780 11296 8832
rect 11336 8780 11388 8832
rect 12348 8780 12400 8832
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 13544 8848 13596 8900
rect 18696 8848 18748 8900
rect 20444 8916 20496 8968
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 23296 9120 23348 9172
rect 22100 9052 22152 9104
rect 20904 8984 20956 9036
rect 22376 8916 22428 8968
rect 22836 9052 22888 9104
rect 24400 9052 24452 9104
rect 23388 8984 23440 9036
rect 23480 8916 23532 8968
rect 25228 8984 25280 9036
rect 22928 8891 22980 8900
rect 22928 8857 22937 8891
rect 22937 8857 22971 8891
rect 22971 8857 22980 8891
rect 22928 8848 22980 8857
rect 13268 8780 13320 8832
rect 19064 8780 19116 8832
rect 21548 8780 21600 8832
rect 25044 8891 25096 8900
rect 25044 8857 25053 8891
rect 25053 8857 25087 8891
rect 25087 8857 25096 8891
rect 25044 8848 25096 8857
rect 25596 8959 25648 8968
rect 25596 8925 25605 8959
rect 25605 8925 25639 8959
rect 25639 8925 25648 8959
rect 25596 8916 25648 8925
rect 25320 8848 25372 8900
rect 24492 8780 24544 8832
rect 25780 8823 25832 8832
rect 25780 8789 25789 8823
rect 25789 8789 25823 8823
rect 25823 8789 25832 8823
rect 25780 8780 25832 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 1952 8551 2004 8560
rect 1952 8517 1961 8551
rect 1961 8517 1995 8551
rect 1995 8517 2004 8551
rect 1952 8508 2004 8517
rect 3056 8508 3108 8560
rect 2780 8372 2832 8424
rect 2964 8440 3016 8492
rect 5816 8576 5868 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 3240 8508 3292 8560
rect 3608 8508 3660 8560
rect 4528 8551 4580 8560
rect 4528 8517 4537 8551
rect 4537 8517 4571 8551
rect 4571 8517 4580 8551
rect 4528 8508 4580 8517
rect 5264 8508 5316 8560
rect 1952 8236 2004 8288
rect 3148 8236 3200 8288
rect 3240 8236 3292 8288
rect 3792 8236 3844 8288
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5632 8440 5684 8492
rect 7380 8508 7432 8560
rect 8760 8576 8812 8628
rect 9036 8576 9088 8628
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 8024 8372 8076 8424
rect 9680 8551 9732 8560
rect 9680 8517 9689 8551
rect 9689 8517 9723 8551
rect 9723 8517 9732 8551
rect 9680 8508 9732 8517
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11520 8576 11572 8628
rect 12716 8576 12768 8628
rect 12072 8508 12124 8560
rect 13820 8576 13872 8628
rect 9312 8440 9364 8492
rect 11612 8440 11664 8492
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11244 8372 11296 8424
rect 9588 8347 9640 8356
rect 9588 8313 9597 8347
rect 9597 8313 9631 8347
rect 9631 8313 9640 8347
rect 9588 8304 9640 8313
rect 10232 8304 10284 8356
rect 4620 8236 4672 8288
rect 5448 8236 5500 8288
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 6460 8236 6512 8288
rect 6828 8236 6880 8288
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 11796 8236 11848 8288
rect 12164 8236 12216 8288
rect 12440 8236 12492 8288
rect 12716 8236 12768 8288
rect 13268 8440 13320 8492
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14188 8508 14240 8560
rect 14740 8508 14792 8560
rect 17592 8508 17644 8560
rect 17868 8508 17920 8560
rect 18420 8508 18472 8560
rect 14096 8483 14148 8492
rect 14096 8449 14130 8483
rect 14130 8449 14148 8483
rect 14096 8440 14148 8449
rect 14556 8440 14608 8492
rect 13636 8372 13688 8424
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 13728 8372 13780 8381
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 16856 8440 16908 8492
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 20260 8576 20312 8628
rect 20720 8576 20772 8628
rect 20996 8576 21048 8628
rect 22192 8576 22244 8628
rect 23020 8576 23072 8628
rect 23388 8576 23440 8628
rect 18696 8551 18748 8560
rect 18696 8517 18705 8551
rect 18705 8517 18739 8551
rect 18739 8517 18748 8551
rect 18696 8508 18748 8517
rect 20904 8508 20956 8560
rect 19064 8483 19116 8492
rect 19064 8449 19073 8483
rect 19073 8449 19107 8483
rect 19107 8449 19116 8483
rect 19064 8440 19116 8449
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 13360 8304 13412 8356
rect 18420 8372 18472 8424
rect 18972 8415 19024 8424
rect 17776 8304 17828 8356
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 21548 8483 21600 8492
rect 21548 8449 21557 8483
rect 21557 8449 21591 8483
rect 21591 8449 21600 8483
rect 21548 8440 21600 8449
rect 22100 8483 22152 8492
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22376 8483 22428 8492
rect 22376 8449 22385 8483
rect 22385 8449 22419 8483
rect 22419 8449 22428 8483
rect 22376 8440 22428 8449
rect 23112 8483 23164 8492
rect 23112 8449 23121 8483
rect 23121 8449 23155 8483
rect 23155 8449 23164 8483
rect 23112 8440 23164 8449
rect 22836 8372 22888 8424
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 23756 8440 23808 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 25596 8440 25648 8492
rect 20996 8304 21048 8356
rect 23480 8304 23532 8356
rect 24860 8304 24912 8356
rect 20720 8236 20772 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2780 8032 2832 8084
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 7380 8032 7432 8084
rect 11520 8032 11572 8084
rect 11796 8032 11848 8084
rect 3332 7964 3384 8016
rect 2596 7760 2648 7812
rect 2320 7692 2372 7744
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5540 7964 5592 8016
rect 6092 7964 6144 8016
rect 5724 7896 5776 7948
rect 5816 7896 5868 7948
rect 11060 7964 11112 8016
rect 10416 7896 10468 7948
rect 10968 7896 11020 7948
rect 11704 7896 11756 7948
rect 12532 7896 12584 7948
rect 4712 7828 4764 7880
rect 3516 7692 3568 7744
rect 4344 7760 4396 7812
rect 5264 7828 5316 7880
rect 5908 7828 5960 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 6644 7871 6696 7880
rect 6644 7837 6654 7871
rect 6654 7837 6688 7871
rect 6688 7837 6696 7871
rect 6644 7828 6696 7837
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7196 7828 7248 7880
rect 10508 7828 10560 7880
rect 6368 7760 6420 7812
rect 4620 7692 4672 7744
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 5816 7735 5868 7744
rect 5816 7701 5825 7735
rect 5825 7701 5859 7735
rect 5859 7701 5868 7735
rect 5816 7692 5868 7701
rect 9128 7760 9180 7812
rect 7104 7692 7156 7744
rect 8024 7692 8076 7744
rect 8760 7735 8812 7744
rect 8760 7701 8769 7735
rect 8769 7701 8803 7735
rect 8803 7701 8812 7735
rect 10968 7760 11020 7812
rect 11244 7828 11296 7880
rect 12624 7828 12676 7880
rect 13268 7896 13320 7948
rect 13452 7896 13504 7948
rect 15200 8032 15252 8084
rect 17408 8075 17460 8084
rect 17408 8041 17417 8075
rect 17417 8041 17451 8075
rect 17451 8041 17460 8075
rect 17408 8032 17460 8041
rect 19248 8032 19300 8084
rect 20904 8032 20956 8084
rect 12072 7760 12124 7812
rect 12348 7803 12400 7812
rect 12348 7769 12357 7803
rect 12357 7769 12391 7803
rect 12391 7769 12400 7803
rect 12348 7760 12400 7769
rect 12532 7760 12584 7812
rect 18052 8007 18104 8016
rect 18052 7973 18061 8007
rect 18061 7973 18095 8007
rect 18095 7973 18104 8007
rect 18052 7964 18104 7973
rect 20628 7964 20680 8016
rect 17040 7896 17092 7948
rect 14188 7828 14240 7880
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 20076 7896 20128 7948
rect 15568 7760 15620 7812
rect 20812 7828 20864 7880
rect 23940 7896 23992 7948
rect 23112 7828 23164 7880
rect 8760 7692 8812 7701
rect 11428 7692 11480 7744
rect 12440 7735 12492 7744
rect 12440 7701 12449 7735
rect 12449 7701 12483 7735
rect 12483 7701 12492 7735
rect 12440 7692 12492 7701
rect 15844 7692 15896 7744
rect 16580 7692 16632 7744
rect 19064 7735 19116 7744
rect 19064 7701 19073 7735
rect 19073 7701 19107 7735
rect 19107 7701 19116 7735
rect 19064 7692 19116 7701
rect 20996 7803 21048 7812
rect 20996 7769 21030 7803
rect 21030 7769 21048 7803
rect 20996 7760 21048 7769
rect 21824 7760 21876 7812
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 23756 7828 23808 7880
rect 24492 7828 24544 7880
rect 24032 7760 24084 7812
rect 21272 7692 21324 7744
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22376 7692 22428 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 25688 7692 25740 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3792 7488 3844 7540
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 4620 7488 4672 7540
rect 6644 7488 6696 7540
rect 3608 7420 3660 7472
rect 5540 7420 5592 7472
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 11612 7488 11664 7540
rect 16580 7488 16632 7540
rect 16764 7488 16816 7540
rect 19064 7488 19116 7540
rect 2320 7395 2372 7404
rect 2320 7361 2354 7395
rect 2354 7361 2372 7395
rect 2320 7352 2372 7361
rect 4620 7352 4672 7404
rect 1952 7284 2004 7336
rect 3424 7284 3476 7336
rect 3240 7148 3292 7200
rect 3516 7148 3568 7200
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7288 7352 7340 7404
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 8116 7352 8168 7404
rect 8484 7352 8536 7404
rect 7932 7216 7984 7268
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10876 7352 10928 7404
rect 12440 7420 12492 7472
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 15568 7420 15620 7472
rect 18696 7420 18748 7472
rect 15384 7395 15436 7404
rect 15384 7361 15418 7395
rect 15418 7361 15436 7395
rect 15384 7352 15436 7361
rect 16856 7395 16908 7404
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 8484 7148 8536 7200
rect 11888 7284 11940 7336
rect 12072 7284 12124 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 13452 7284 13504 7336
rect 11336 7259 11388 7268
rect 11336 7225 11345 7259
rect 11345 7225 11379 7259
rect 11379 7225 11388 7259
rect 11336 7216 11388 7225
rect 11612 7259 11664 7268
rect 11612 7225 11621 7259
rect 11621 7225 11655 7259
rect 11655 7225 11664 7259
rect 11612 7216 11664 7225
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 19432 7352 19484 7404
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 20996 7488 21048 7540
rect 20444 7420 20496 7472
rect 19984 7216 20036 7268
rect 11980 7191 12032 7200
rect 11980 7157 11989 7191
rect 11989 7157 12023 7191
rect 12023 7157 12032 7191
rect 11980 7148 12032 7157
rect 16948 7148 17000 7200
rect 19340 7148 19392 7200
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 20812 7352 20864 7404
rect 22008 7488 22060 7540
rect 21824 7463 21876 7472
rect 21824 7429 21833 7463
rect 21833 7429 21867 7463
rect 21867 7429 21876 7463
rect 21824 7420 21876 7429
rect 23296 7420 23348 7472
rect 24308 7488 24360 7540
rect 25044 7488 25096 7540
rect 25596 7488 25648 7540
rect 26148 7488 26200 7540
rect 20996 7284 21048 7336
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 22468 7284 22520 7336
rect 22652 7327 22704 7336
rect 22652 7293 22661 7327
rect 22661 7293 22695 7327
rect 22695 7293 22704 7327
rect 22652 7284 22704 7293
rect 22192 7216 22244 7268
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 23848 7420 23900 7472
rect 23940 7395 23992 7404
rect 23940 7361 23949 7395
rect 23949 7361 23983 7395
rect 23983 7361 23992 7395
rect 23940 7352 23992 7361
rect 24032 7352 24084 7404
rect 24676 7352 24728 7404
rect 25688 7352 25740 7404
rect 23480 7216 23532 7268
rect 20628 7148 20680 7200
rect 20904 7148 20956 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 7840 6944 7892 6996
rect 1952 6851 2004 6860
rect 1952 6817 1961 6851
rect 1961 6817 1995 6851
rect 1995 6817 2004 6851
rect 1952 6808 2004 6817
rect 3608 6808 3660 6860
rect 11428 6944 11480 6996
rect 11980 6944 12032 6996
rect 12624 6944 12676 6996
rect 14280 6944 14332 6996
rect 16120 6944 16172 6996
rect 19156 6944 19208 6996
rect 3240 6740 3292 6792
rect 3884 6740 3936 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4620 6740 4672 6792
rect 5816 6740 5868 6792
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 11060 6876 11112 6928
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 2320 6672 2372 6724
rect 3148 6672 3200 6724
rect 2136 6604 2188 6656
rect 3700 6604 3752 6656
rect 8852 6672 8904 6724
rect 10508 6672 10560 6724
rect 11336 6783 11388 6792
rect 11336 6749 11370 6783
rect 11370 6749 11388 6783
rect 11336 6740 11388 6749
rect 13820 6740 13872 6792
rect 14648 6740 14700 6792
rect 16856 6808 16908 6860
rect 18604 6876 18656 6928
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 11888 6672 11940 6724
rect 14280 6715 14332 6724
rect 14280 6681 14289 6715
rect 14289 6681 14323 6715
rect 14323 6681 14332 6715
rect 14280 6672 14332 6681
rect 4620 6604 4672 6656
rect 7748 6604 7800 6656
rect 8116 6604 8168 6656
rect 11336 6604 11388 6656
rect 14556 6604 14608 6656
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 18052 6740 18104 6792
rect 18880 6808 18932 6860
rect 19432 6944 19484 6996
rect 21548 6944 21600 6996
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 18696 6783 18748 6792
rect 18696 6749 18705 6783
rect 18705 6749 18739 6783
rect 18739 6749 18748 6783
rect 18696 6740 18748 6749
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19156 6740 19208 6792
rect 21456 6808 21508 6860
rect 24216 6944 24268 6996
rect 24584 6944 24636 6996
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 20996 6783 21048 6792
rect 20996 6749 21005 6783
rect 21005 6749 21039 6783
rect 21039 6749 21048 6783
rect 20996 6740 21048 6749
rect 15568 6672 15620 6724
rect 16856 6672 16908 6724
rect 15936 6604 15988 6656
rect 16028 6604 16080 6656
rect 17960 6604 18012 6656
rect 18972 6672 19024 6724
rect 21272 6740 21324 6792
rect 22468 6808 22520 6860
rect 23480 6851 23532 6860
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23480 6808 23532 6817
rect 22928 6740 22980 6792
rect 24676 6876 24728 6928
rect 21732 6672 21784 6724
rect 22100 6672 22152 6724
rect 20720 6604 20772 6656
rect 21364 6647 21416 6656
rect 21364 6613 21373 6647
rect 21373 6613 21407 6647
rect 21407 6613 21416 6647
rect 21364 6604 21416 6613
rect 23020 6715 23072 6724
rect 23020 6681 23029 6715
rect 23029 6681 23063 6715
rect 23063 6681 23072 6715
rect 23020 6672 23072 6681
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 24952 6783 25004 6792
rect 24952 6749 24961 6783
rect 24961 6749 24995 6783
rect 24995 6749 25004 6783
rect 24952 6740 25004 6749
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 24768 6715 24820 6724
rect 24768 6681 24777 6715
rect 24777 6681 24811 6715
rect 24811 6681 24820 6715
rect 24768 6672 24820 6681
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 25412 6647 25464 6656
rect 25412 6613 25421 6647
rect 25421 6613 25455 6647
rect 25455 6613 25464 6647
rect 25412 6604 25464 6613
rect 25780 6647 25832 6656
rect 25780 6613 25789 6647
rect 25789 6613 25823 6647
rect 25823 6613 25832 6647
rect 25780 6604 25832 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2136 6375 2188 6384
rect 2136 6341 2145 6375
rect 2145 6341 2179 6375
rect 2179 6341 2188 6375
rect 2136 6332 2188 6341
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 4068 6400 4120 6452
rect 6460 6400 6512 6452
rect 6552 6400 6604 6452
rect 8116 6443 8168 6452
rect 8116 6409 8125 6443
rect 8125 6409 8159 6443
rect 8159 6409 8168 6443
rect 8116 6400 8168 6409
rect 8852 6400 8904 6452
rect 2596 6264 2648 6316
rect 4620 6332 4672 6384
rect 5264 6332 5316 6384
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 6460 6264 6512 6316
rect 7932 6332 7984 6384
rect 8300 6332 8352 6384
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8392 6264 8444 6316
rect 8484 6264 8536 6316
rect 8944 6264 8996 6316
rect 9312 6264 9364 6316
rect 10968 6400 11020 6452
rect 14188 6400 14240 6452
rect 15384 6400 15436 6452
rect 15936 6400 15988 6452
rect 12072 6332 12124 6384
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 14096 6264 14148 6316
rect 15476 6332 15528 6384
rect 24400 6400 24452 6452
rect 19340 6375 19392 6384
rect 19340 6341 19374 6375
rect 19374 6341 19392 6375
rect 19340 6332 19392 6341
rect 15568 6264 15620 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 15936 6307 15988 6316
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 16028 6307 16080 6316
rect 16028 6273 16037 6307
rect 16037 6273 16071 6307
rect 16071 6273 16080 6307
rect 16028 6264 16080 6273
rect 11336 6239 11388 6248
rect 11336 6205 11345 6239
rect 11345 6205 11379 6239
rect 11379 6205 11388 6239
rect 11336 6196 11388 6205
rect 11980 6196 12032 6248
rect 14740 6196 14792 6248
rect 16764 6264 16816 6316
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 19800 6264 19852 6316
rect 21272 6307 21324 6316
rect 21272 6273 21281 6307
rect 21281 6273 21315 6307
rect 21315 6273 21324 6307
rect 21272 6264 21324 6273
rect 16396 6196 16448 6248
rect 3424 6128 3476 6180
rect 4160 6128 4212 6180
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 2596 6060 2648 6112
rect 8392 6128 8444 6180
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5724 6060 5776 6112
rect 8300 6060 8352 6112
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 14464 6128 14516 6180
rect 16212 6128 16264 6180
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 20260 6196 20312 6248
rect 21456 6264 21508 6316
rect 21732 6264 21784 6316
rect 23020 6264 23072 6316
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 23296 6307 23348 6316
rect 23296 6273 23305 6307
rect 23305 6273 23339 6307
rect 23339 6273 23348 6307
rect 23296 6264 23348 6273
rect 25596 6332 25648 6384
rect 23756 6264 23808 6316
rect 24676 6264 24728 6316
rect 22560 6196 22612 6248
rect 22652 6196 22704 6248
rect 24768 6196 24820 6248
rect 20536 6128 20588 6180
rect 21732 6128 21784 6180
rect 24952 6128 25004 6180
rect 10784 6060 10836 6112
rect 13912 6060 13964 6112
rect 14280 6060 14332 6112
rect 15936 6060 15988 6112
rect 17408 6060 17460 6112
rect 19800 6060 19852 6112
rect 20904 6060 20956 6112
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 24032 6060 24084 6112
rect 25136 6103 25188 6112
rect 25136 6069 25145 6103
rect 25145 6069 25179 6103
rect 25179 6069 25188 6103
rect 25136 6060 25188 6069
rect 25320 6128 25372 6180
rect 25596 6060 25648 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2504 5856 2556 5908
rect 4436 5856 4488 5908
rect 5264 5856 5316 5908
rect 5540 5856 5592 5908
rect 6552 5788 6604 5840
rect 2688 5652 2740 5704
rect 3148 5652 3200 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 2596 5584 2648 5636
rect 6092 5652 6144 5704
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 15292 5856 15344 5908
rect 15844 5856 15896 5908
rect 18328 5856 18380 5908
rect 21732 5856 21784 5908
rect 22100 5856 22152 5908
rect 23112 5856 23164 5908
rect 23940 5856 23992 5908
rect 25320 5856 25372 5908
rect 25780 5899 25832 5908
rect 25780 5865 25789 5899
rect 25789 5865 25823 5899
rect 25823 5865 25832 5899
rect 25780 5856 25832 5865
rect 8300 5788 8352 5840
rect 13820 5788 13872 5840
rect 14188 5788 14240 5840
rect 14740 5788 14792 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 17224 5788 17276 5840
rect 17684 5831 17736 5840
rect 17684 5797 17693 5831
rect 17693 5797 17727 5831
rect 17727 5797 17736 5831
rect 17684 5788 17736 5797
rect 19340 5788 19392 5840
rect 20536 5788 20588 5840
rect 23756 5788 23808 5840
rect 8760 5720 8812 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 10784 5695 10836 5704
rect 10784 5661 10818 5695
rect 10818 5661 10836 5695
rect 10784 5652 10836 5661
rect 14004 5720 14056 5772
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 5540 5627 5592 5636
rect 5540 5593 5574 5627
rect 5574 5593 5592 5627
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 5540 5584 5592 5593
rect 7748 5584 7800 5636
rect 9312 5584 9364 5636
rect 9496 5584 9548 5636
rect 13820 5584 13872 5636
rect 14096 5584 14148 5636
rect 6460 5516 6512 5568
rect 6644 5516 6696 5568
rect 8668 5516 8720 5568
rect 11980 5516 12032 5568
rect 14556 5516 14608 5568
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 16764 5720 16816 5772
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 15660 5652 15712 5704
rect 17776 5720 17828 5772
rect 19064 5720 19116 5772
rect 15844 5627 15896 5636
rect 15844 5593 15878 5627
rect 15878 5593 15896 5627
rect 15844 5584 15896 5593
rect 17224 5627 17276 5636
rect 17224 5593 17233 5627
rect 17233 5593 17267 5627
rect 17267 5593 17276 5627
rect 17224 5584 17276 5593
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 22192 5652 22244 5704
rect 22652 5652 22704 5704
rect 16120 5516 16172 5568
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 20812 5584 20864 5636
rect 21364 5584 21416 5636
rect 21548 5584 21600 5636
rect 23940 5584 23992 5636
rect 24032 5627 24084 5636
rect 24032 5593 24041 5627
rect 24041 5593 24075 5627
rect 24075 5593 24084 5627
rect 24032 5584 24084 5593
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24860 5652 24912 5704
rect 24768 5627 24820 5636
rect 24768 5593 24777 5627
rect 24777 5593 24811 5627
rect 24811 5593 24820 5627
rect 24768 5584 24820 5593
rect 25596 5695 25648 5704
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 25504 5584 25556 5636
rect 21272 5516 21324 5568
rect 22100 5559 22152 5568
rect 22100 5525 22109 5559
rect 22109 5525 22143 5559
rect 22143 5525 22152 5559
rect 22100 5516 22152 5525
rect 23296 5516 23348 5568
rect 23480 5516 23532 5568
rect 23664 5516 23716 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1952 5312 2004 5364
rect 3240 5312 3292 5364
rect 5540 5355 5592 5364
rect 5540 5321 5549 5355
rect 5549 5321 5583 5355
rect 5583 5321 5592 5355
rect 5540 5312 5592 5321
rect 5816 5312 5868 5364
rect 6092 5312 6144 5364
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 4620 5287 4672 5296
rect 4620 5253 4629 5287
rect 4629 5253 4663 5287
rect 4663 5253 4672 5287
rect 4620 5244 4672 5253
rect 6460 5244 6512 5296
rect 8576 5312 8628 5364
rect 7472 5287 7524 5296
rect 5264 5176 5316 5228
rect 7472 5253 7481 5287
rect 7481 5253 7515 5287
rect 7515 5253 7524 5287
rect 7472 5244 7524 5253
rect 7932 5244 7984 5296
rect 8760 5244 8812 5296
rect 8668 5176 8720 5228
rect 13176 5176 13228 5228
rect 14464 5312 14516 5364
rect 15844 5312 15896 5364
rect 19432 5312 19484 5364
rect 14648 5244 14700 5296
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2504 5040 2556 5092
rect 2596 5040 2648 5092
rect 4620 5040 4672 5092
rect 7932 5083 7984 5092
rect 7932 5049 7941 5083
rect 7941 5049 7975 5083
rect 7975 5049 7984 5083
rect 7932 5040 7984 5049
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 6644 4972 6696 5024
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 14096 5176 14148 5228
rect 15108 5176 15160 5228
rect 14648 5108 14700 5160
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 14188 5040 14240 5092
rect 15384 4972 15436 5024
rect 15752 5176 15804 5228
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 17040 5244 17092 5296
rect 18236 5244 18288 5296
rect 15844 5108 15896 5160
rect 16396 5219 16448 5228
rect 16396 5185 16405 5219
rect 16405 5185 16439 5219
rect 16439 5185 16448 5219
rect 16396 5176 16448 5185
rect 18052 5176 18104 5228
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 20260 5219 20312 5228
rect 20260 5185 20269 5219
rect 20269 5185 20303 5219
rect 20303 5185 20312 5219
rect 20260 5176 20312 5185
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 20996 5312 21048 5364
rect 21272 5312 21324 5364
rect 20812 5244 20864 5296
rect 22100 5312 22152 5364
rect 20444 5176 20496 5228
rect 21272 5219 21324 5228
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 21456 5219 21508 5228
rect 21456 5185 21465 5219
rect 21465 5185 21499 5219
rect 21499 5185 21508 5219
rect 21456 5176 21508 5185
rect 21732 5176 21784 5228
rect 22192 5244 22244 5296
rect 23296 5244 23348 5296
rect 25320 5312 25372 5364
rect 23020 5176 23072 5228
rect 23480 5176 23532 5228
rect 23204 5108 23256 5160
rect 23848 5176 23900 5228
rect 25780 5355 25832 5364
rect 25780 5321 25789 5355
rect 25789 5321 25823 5355
rect 25823 5321 25832 5355
rect 25780 5312 25832 5321
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20536 5040 20588 5092
rect 23664 5040 23716 5092
rect 23848 5040 23900 5092
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2780 4768 2832 4820
rect 8392 4768 8444 4820
rect 13820 4768 13872 4820
rect 14648 4768 14700 4820
rect 14740 4768 14792 4820
rect 15476 4768 15528 4820
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18880 4811 18932 4820
rect 18880 4777 18889 4811
rect 18889 4777 18923 4811
rect 18923 4777 18932 4811
rect 18880 4768 18932 4777
rect 1952 4632 2004 4684
rect 2228 4564 2280 4616
rect 8484 4632 8536 4684
rect 16764 4632 16816 4684
rect 8300 4564 8352 4616
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13268 4564 13320 4616
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 17960 4564 18012 4616
rect 18328 4700 18380 4752
rect 20996 4768 21048 4820
rect 21456 4768 21508 4820
rect 21732 4768 21784 4820
rect 25504 4768 25556 4820
rect 12808 4428 12860 4480
rect 14004 4428 14056 4480
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 16120 4539 16172 4548
rect 16120 4505 16129 4539
rect 16129 4505 16163 4539
rect 16163 4505 16172 4539
rect 16120 4496 16172 4505
rect 16212 4539 16264 4548
rect 16212 4505 16221 4539
rect 16221 4505 16255 4539
rect 16255 4505 16264 4539
rect 16212 4496 16264 4505
rect 17684 4496 17736 4548
rect 18880 4564 18932 4616
rect 18972 4564 19024 4616
rect 21824 4700 21876 4752
rect 19432 4607 19484 4616
rect 19432 4573 19441 4607
rect 19441 4573 19475 4607
rect 19475 4573 19484 4607
rect 19432 4564 19484 4573
rect 20260 4564 20312 4616
rect 23204 4632 23256 4684
rect 23296 4632 23348 4684
rect 21640 4564 21692 4616
rect 23020 4564 23072 4616
rect 17040 4428 17092 4480
rect 19524 4496 19576 4548
rect 21548 4496 21600 4548
rect 19432 4428 19484 4480
rect 21732 4428 21784 4480
rect 23756 4607 23808 4616
rect 23756 4573 23765 4607
rect 23765 4573 23799 4607
rect 23799 4573 23808 4607
rect 23756 4564 23808 4573
rect 23848 4607 23900 4616
rect 23848 4573 23857 4607
rect 23857 4573 23891 4607
rect 23891 4573 23900 4607
rect 23848 4564 23900 4573
rect 24124 4564 24176 4616
rect 23296 4496 23348 4548
rect 23112 4428 23164 4480
rect 24860 4496 24912 4548
rect 24768 4428 24820 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 14740 4224 14792 4276
rect 17408 4224 17460 4276
rect 19616 4267 19668 4276
rect 19616 4233 19625 4267
rect 19625 4233 19659 4267
rect 19659 4233 19668 4267
rect 19616 4224 19668 4233
rect 20168 4224 20220 4276
rect 14096 4088 14148 4140
rect 14372 4088 14424 4140
rect 12532 4020 12584 4072
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 15292 4020 15344 4072
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 15844 4088 15896 4140
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 15936 4020 15988 4072
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 16396 4131 16448 4140
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 16764 4156 16816 4208
rect 18880 4156 18932 4208
rect 19800 4156 19852 4208
rect 16948 4088 17000 4140
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 17500 4131 17552 4140
rect 17500 4097 17509 4131
rect 17509 4097 17543 4131
rect 17543 4097 17552 4131
rect 17500 4088 17552 4097
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 19248 4088 19300 4140
rect 13728 3884 13780 3936
rect 13820 3884 13872 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15660 3952 15712 4004
rect 16580 3952 16632 4004
rect 17684 4020 17736 4072
rect 16488 3884 16540 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 19432 4020 19484 4072
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20536 4199 20588 4208
rect 20536 4165 20545 4199
rect 20545 4165 20579 4199
rect 20579 4165 20588 4199
rect 20536 4156 20588 4165
rect 21548 4224 21600 4276
rect 22100 4224 22152 4276
rect 22560 4224 22612 4276
rect 23020 4224 23072 4276
rect 23112 4224 23164 4276
rect 19708 3952 19760 4004
rect 20444 4088 20496 4140
rect 21456 4199 21508 4208
rect 21456 4165 21465 4199
rect 21465 4165 21499 4199
rect 21499 4165 21508 4199
rect 21456 4156 21508 4165
rect 20536 4020 20588 4072
rect 21364 4088 21416 4140
rect 21732 4088 21784 4140
rect 20444 3952 20496 4004
rect 22100 4131 22152 4140
rect 22100 4097 22109 4131
rect 22109 4097 22143 4131
rect 22143 4097 22152 4131
rect 22100 4088 22152 4097
rect 22836 4088 22888 4140
rect 23020 4131 23072 4140
rect 23020 4097 23029 4131
rect 23029 4097 23063 4131
rect 23063 4097 23072 4131
rect 23020 4088 23072 4097
rect 23572 4156 23624 4208
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 22284 4020 22336 4072
rect 24768 4088 24820 4140
rect 24860 4131 24912 4140
rect 24860 4097 24869 4131
rect 24869 4097 24903 4131
rect 24903 4097 24912 4131
rect 24860 4088 24912 4097
rect 25504 4088 25556 4140
rect 25412 3995 25464 4004
rect 25412 3961 25421 3995
rect 25421 3961 25455 3995
rect 25455 3961 25464 3995
rect 25412 3952 25464 3961
rect 25780 3995 25832 4004
rect 25780 3961 25789 3995
rect 25789 3961 25823 3995
rect 25823 3961 25832 3995
rect 25780 3952 25832 3961
rect 21180 3884 21232 3936
rect 22468 3927 22520 3936
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 22468 3884 22520 3893
rect 22928 3884 22980 3936
rect 23112 3884 23164 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 16120 3680 16172 3732
rect 16488 3680 16540 3732
rect 18972 3723 19024 3732
rect 18972 3689 18981 3723
rect 18981 3689 19015 3723
rect 19015 3689 19024 3723
rect 18972 3680 19024 3689
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 18696 3655 18748 3664
rect 18696 3621 18705 3655
rect 18705 3621 18739 3655
rect 18739 3621 18748 3655
rect 18696 3612 18748 3621
rect 19340 3544 19392 3596
rect 19432 3544 19484 3596
rect 13728 3476 13780 3528
rect 15476 3476 15528 3528
rect 18144 3476 18196 3528
rect 19800 3544 19852 3596
rect 23112 3680 23164 3732
rect 23572 3680 23624 3732
rect 24768 3680 24820 3732
rect 23388 3612 23440 3664
rect 19708 3519 19760 3528
rect 19708 3485 19717 3519
rect 19717 3485 19751 3519
rect 19751 3485 19760 3519
rect 19708 3476 19760 3485
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 23480 3544 23532 3596
rect 14372 3451 14424 3460
rect 14372 3417 14406 3451
rect 14406 3417 14424 3451
rect 14372 3408 14424 3417
rect 16672 3408 16724 3460
rect 17776 3408 17828 3460
rect 18788 3408 18840 3460
rect 19340 3408 19392 3460
rect 20536 3476 20588 3528
rect 16948 3340 17000 3392
rect 17684 3340 17736 3392
rect 19432 3340 19484 3392
rect 20260 3340 20312 3392
rect 20352 3340 20404 3392
rect 21180 3340 21232 3392
rect 21548 3476 21600 3528
rect 22468 3519 22520 3528
rect 21824 3451 21876 3460
rect 21824 3417 21842 3451
rect 21842 3417 21876 3451
rect 21824 3408 21876 3417
rect 22468 3485 22502 3519
rect 22502 3485 22520 3519
rect 22468 3476 22520 3485
rect 24124 3476 24176 3528
rect 23480 3408 23532 3460
rect 22836 3340 22888 3392
rect 23020 3340 23072 3392
rect 23848 3451 23900 3460
rect 23848 3417 23857 3451
rect 23857 3417 23891 3451
rect 23891 3417 23900 3451
rect 23848 3408 23900 3417
rect 24492 3476 24544 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 25780 3383 25832 3392
rect 25780 3349 25789 3383
rect 25789 3349 25823 3383
rect 25823 3349 25832 3383
rect 25780 3340 25832 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 15568 3136 15620 3188
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 16764 3136 16816 3188
rect 15108 3068 15160 3120
rect 15292 3068 15344 3120
rect 16120 3068 16172 3120
rect 16580 3068 16632 3120
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 15200 2864 15252 2916
rect 15936 2932 15988 2984
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17316 3136 17368 3188
rect 18328 3068 18380 3120
rect 18696 3068 18748 3120
rect 19616 3136 19668 3188
rect 19800 3179 19852 3188
rect 19800 3145 19809 3179
rect 19809 3145 19843 3179
rect 19843 3145 19852 3179
rect 19800 3136 19852 3145
rect 19892 3136 19944 3188
rect 20352 3136 20404 3188
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 17408 3000 17460 3052
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 17040 2864 17092 2916
rect 17316 2864 17368 2916
rect 18788 3000 18840 3052
rect 19524 3000 19576 3052
rect 19708 3000 19760 3052
rect 20260 3000 20312 3052
rect 20628 3111 20680 3120
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 21088 3136 21140 3188
rect 21824 3179 21876 3188
rect 21824 3145 21833 3179
rect 21833 3145 21867 3179
rect 21867 3145 21876 3179
rect 21824 3136 21876 3145
rect 20996 3068 21048 3120
rect 22192 3136 22244 3188
rect 22468 3136 22520 3188
rect 23296 3136 23348 3188
rect 23848 3136 23900 3188
rect 24492 3179 24544 3188
rect 24492 3145 24501 3179
rect 24501 3145 24535 3179
rect 24535 3145 24544 3179
rect 24492 3136 24544 3145
rect 22928 3111 22980 3120
rect 20168 2932 20220 2984
rect 20904 3043 20956 3052
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 21088 3043 21140 3052
rect 21088 3009 21097 3043
rect 21097 3009 21131 3043
rect 21131 3009 21140 3043
rect 21088 3000 21140 3009
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 21364 3000 21416 3052
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 22468 3043 22520 3052
rect 22468 3009 22477 3043
rect 22477 3009 22511 3043
rect 22511 3009 22520 3043
rect 22468 3000 22520 3009
rect 22928 3077 22962 3111
rect 22962 3077 22980 3111
rect 22928 3068 22980 3077
rect 23112 3068 23164 3120
rect 24124 3111 24176 3120
rect 24124 3077 24133 3111
rect 24133 3077 24167 3111
rect 24167 3077 24176 3111
rect 24124 3068 24176 3077
rect 24860 3000 24912 3052
rect 25228 3000 25280 3052
rect 22560 2932 22612 2984
rect 18604 2796 18656 2848
rect 19340 2796 19392 2848
rect 19892 2796 19944 2848
rect 20536 2796 20588 2848
rect 20996 2796 21048 2848
rect 21088 2796 21140 2848
rect 21548 2796 21600 2848
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10416 2592 10468 2644
rect 18604 2592 18656 2644
rect 18696 2524 18748 2576
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 17960 2456 18012 2508
rect 10324 2388 10376 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12256 2388 12308 2440
rect 13820 2388 13872 2440
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14004 2388 14056 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16120 2388 16172 2440
rect 16856 2388 16908 2440
rect 17224 2388 17276 2440
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19432 2456 19484 2508
rect 21272 2592 21324 2644
rect 20352 2524 20404 2576
rect 22284 2524 22336 2576
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 20904 2456 20956 2508
rect 19708 2388 19760 2440
rect 20444 2388 20496 2440
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 21088 2388 21140 2440
rect 21916 2388 21968 2440
rect 20076 2320 20128 2372
rect 23020 2388 23072 2440
rect 23204 2388 23256 2440
rect 23848 2388 23900 2440
rect 24860 2431 24912 2440
rect 24860 2397 24869 2431
rect 24869 2397 24903 2431
rect 24903 2397 24912 2431
rect 24860 2388 24912 2397
rect 11612 2252 11664 2304
rect 12900 2252 12952 2304
rect 13544 2252 13596 2304
rect 14188 2252 14240 2304
rect 14832 2252 14884 2304
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 16764 2252 16816 2304
rect 17408 2252 17460 2304
rect 18052 2252 18104 2304
rect 19432 2252 19484 2304
rect 19984 2252 20036 2304
rect 20628 2252 20680 2304
rect 21180 2252 21232 2304
rect 22560 2252 22612 2304
rect 23204 2252 23256 2304
rect 23848 2252 23900 2304
rect 24492 2252 24544 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 12898 28676 12954 29476
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 12912 27130 12940 28676
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 110 25664 166 25673
rect 110 25599 166 25608
rect 124 14074 152 25599
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 9416 23866 9444 24754
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 10888 23730 10916 24618
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10980 23730 11008 24006
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 4620 23588 4672 23594
rect 4620 23530 4672 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3608 23248 3660 23254
rect 3608 23190 3660 23196
rect 3700 23248 3752 23254
rect 4632 23202 4660 23530
rect 3700 23190 3752 23196
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1964 22506 1992 23054
rect 2504 23044 2556 23050
rect 2504 22986 2556 22992
rect 2516 22778 2544 22986
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2608 22778 2636 22918
rect 3252 22794 3280 23122
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 3160 22766 3280 22794
rect 1952 22500 2004 22506
rect 1952 22442 2004 22448
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 860 21321 888 21490
rect 1964 21486 1992 22442
rect 2504 22094 2556 22098
rect 2608 22094 2636 22714
rect 3160 22574 3188 22766
rect 3620 22642 3648 23190
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 2792 22166 2820 22510
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2504 22092 2636 22094
rect 2556 22066 2636 22092
rect 2504 22034 2556 22040
rect 2412 22024 2464 22030
rect 2332 21984 2412 22012
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2148 21622 2176 21830
rect 2136 21616 2188 21622
rect 2136 21558 2188 21564
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 846 21312 902 21321
rect 846 21247 902 21256
rect 1964 20942 1992 21422
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 2136 20868 2188 20874
rect 2136 20810 2188 20816
rect 2148 20602 2176 20810
rect 2332 20602 2360 21984
rect 2412 21966 2464 21972
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2424 20602 2452 20878
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2412 20596 2464 20602
rect 2412 20538 2464 20544
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 1964 20058 1992 20402
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2240 19718 2268 20198
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19378 2268 19654
rect 2332 19446 2360 20538
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 848 18760 900 18766
rect 848 18702 900 18708
rect 860 18601 888 18702
rect 1952 18624 2004 18630
rect 846 18592 902 18601
rect 1952 18566 2004 18572
rect 846 18527 902 18536
rect 1964 17610 1992 18566
rect 2240 18426 2268 19314
rect 2332 18766 2360 19382
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2424 18290 2452 20538
rect 2516 20466 2544 22034
rect 3160 22030 3188 22510
rect 3620 22438 3648 22578
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3620 22234 3648 22374
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3712 22166 3740 23190
rect 4448 23186 4660 23202
rect 5184 23202 5212 23598
rect 5276 23322 5304 23598
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 4436 23180 4660 23186
rect 4488 23174 4660 23180
rect 4712 23180 4764 23186
rect 4436 23122 4488 23128
rect 4712 23122 4764 23128
rect 5184 23174 5304 23202
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22574 4660 22986
rect 3792 22568 3844 22574
rect 3792 22510 3844 22516
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 3804 22166 3832 22510
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 3700 22160 3752 22166
rect 3700 22102 3752 22108
rect 3792 22160 3844 22166
rect 4540 22137 4568 22170
rect 3792 22102 3844 22108
rect 4526 22128 4582 22137
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 2700 20466 2728 21966
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3620 21690 3648 21898
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3804 21554 3832 22102
rect 4526 22063 4582 22072
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3252 21010 3280 21286
rect 3344 21146 3372 21490
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3436 20942 3464 21286
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 3424 20936 3476 20942
rect 3424 20878 3476 20884
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2516 18834 2544 20402
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 18834 2636 19110
rect 2700 18902 2728 20402
rect 2792 19854 2820 20470
rect 2884 20330 2912 20878
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3252 20534 3280 20742
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 3252 20058 3280 20470
rect 3436 20398 3464 20878
rect 3804 20534 3832 21490
rect 4540 21434 4568 22063
rect 4632 22030 4660 22374
rect 4724 22234 4752 23122
rect 5184 23050 5212 23174
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 4896 22976 4948 22982
rect 4816 22936 4896 22964
rect 4816 22710 4844 22936
rect 4896 22918 4948 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22778 5304 23174
rect 4988 22772 5040 22778
rect 4908 22732 4988 22760
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4908 22438 4936 22732
rect 4988 22714 5040 22720
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4908 22030 4936 22374
rect 5172 22160 5224 22166
rect 5078 22128 5134 22137
rect 5172 22102 5224 22108
rect 5078 22063 5134 22072
rect 5092 22030 5120 22063
rect 5184 22030 5212 22102
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5368 21894 5396 22374
rect 5460 22234 5488 23462
rect 5552 23118 5580 23462
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 6012 22098 6040 23598
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8300 23112 8352 23118
rect 8300 23054 8352 23060
rect 7012 23044 7064 23050
rect 7012 22986 7064 22992
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6380 22166 6408 22918
rect 6656 22710 6684 22918
rect 7024 22778 7052 22986
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 6368 22160 6420 22166
rect 6368 22102 6420 22108
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 6380 22030 6408 22102
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 5920 21894 5948 21966
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4540 21406 4660 21434
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20936 4120 20942
rect 4632 20890 4660 21406
rect 5368 21146 5396 21830
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 4068 20878 4120 20884
rect 4080 20534 4108 20878
rect 4540 20862 4660 20890
rect 4804 20868 4856 20874
rect 3792 20528 3844 20534
rect 3792 20470 3844 20476
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3252 19854 3280 19994
rect 3620 19922 3648 20402
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 2792 19310 2820 19790
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2688 18896 2740 18902
rect 2688 18838 2740 18844
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2792 18698 2820 19246
rect 3160 18834 3188 19382
rect 3804 19378 3832 19994
rect 4080 19922 4108 20470
rect 4540 20466 4568 20862
rect 4804 20810 4856 20816
rect 4620 20800 4672 20806
rect 4620 20742 4672 20748
rect 4632 20466 4660 20742
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3896 19310 3924 19790
rect 4080 19378 4108 19858
rect 4632 19854 4660 20402
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4724 19496 4752 20402
rect 4632 19468 4752 19496
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4632 19310 4660 19468
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2424 18170 2452 18226
rect 2332 18142 2452 18170
rect 2332 17678 2360 18142
rect 2792 17882 2820 18634
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2884 18272 2912 18566
rect 2964 18284 3016 18290
rect 2884 18244 2964 18272
rect 2964 18226 3016 18232
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16250 1624 16390
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1768 16176 1820 16182
rect 1768 16118 1820 16124
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15881 888 16050
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1780 15706 1808 16118
rect 2332 16114 2360 17614
rect 3804 17338 3832 18702
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3804 17202 3832 17274
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3896 17134 3924 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4080 18426 4108 18702
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 4068 18284 4120 18290
rect 4172 18272 4200 18906
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4448 18290 4476 18566
rect 4120 18244 4200 18272
rect 4436 18284 4488 18290
rect 4068 18226 4120 18232
rect 4436 18226 4488 18232
rect 3988 17882 4016 18226
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3988 17678 4016 17818
rect 4080 17796 4108 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4160 17808 4212 17814
rect 4080 17768 4160 17796
rect 4160 17750 4212 17756
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4172 17610 4200 17750
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4448 17202 4476 17478
rect 4632 17338 4660 19246
rect 4724 18766 4752 19314
rect 4816 19281 4844 20810
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5092 19854 5120 20334
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5184 19854 5212 20198
rect 5644 19854 5672 20742
rect 5736 19854 5764 21014
rect 5828 20942 5856 21014
rect 6380 21010 6408 21966
rect 6656 21350 6684 22646
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 6840 21894 6868 22510
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 21706 6868 21830
rect 6840 21690 6960 21706
rect 6840 21684 6972 21690
rect 6840 21678 6920 21684
rect 6920 21626 6972 21632
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6472 21010 6500 21286
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 6000 20936 6052 20942
rect 6052 20896 6316 20924
rect 6000 20878 6052 20884
rect 6288 20890 6316 20896
rect 6472 20890 6500 20946
rect 6288 20862 6500 20890
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4802 19272 4858 19281
rect 4802 19207 4858 19216
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 18766 4844 19110
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5092 18766 5120 18906
rect 5644 18834 5672 19654
rect 5828 19446 5856 19654
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5920 19378 5948 19654
rect 6564 19496 6592 20878
rect 6380 19468 6592 19496
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6012 19258 6040 19314
rect 5920 19230 6040 19258
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 5080 18760 5132 18766
rect 5356 18760 5408 18766
rect 5132 18720 5304 18748
rect 5080 18702 5132 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18426 5304 18720
rect 5356 18702 5408 18708
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5368 17882 5396 18702
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5552 18426 5580 18634
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5736 18358 5764 18770
rect 5816 18760 5868 18766
rect 5920 18748 5948 19230
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 5868 18720 5948 18748
rect 5816 18702 5868 18708
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 5828 18170 5856 18702
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5920 18290 5948 18566
rect 6012 18290 6040 19110
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5828 18142 5948 18170
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16114 3924 17070
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16250 4660 17274
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 2424 15706 2452 16050
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 1504 15065 1532 15370
rect 1490 15056 1546 15065
rect 2608 15026 2636 15642
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 1490 14991 1546 15000
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 112 14068 164 14074
rect 112 14010 164 14016
rect 1596 13938 1624 14350
rect 1872 13938 1900 14758
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 2148 13530 2176 14282
rect 2608 13530 2636 14962
rect 2700 14890 2728 15370
rect 2884 15026 2912 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2608 12442 2636 13466
rect 2700 13258 2728 14826
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 13870 2912 14758
rect 2976 13938 3004 15302
rect 3160 15162 3188 15302
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3068 14414 3096 14894
rect 3160 14482 3188 14962
rect 3252 14618 3280 15506
rect 3344 15434 3372 15506
rect 4080 15502 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 4068 15496 4120 15502
rect 4120 15444 4200 15450
rect 4068 15438 4200 15444
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3344 14822 3372 15370
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3620 14770 3648 15438
rect 3976 15428 4028 15434
rect 4080 15422 4200 15438
rect 3976 15370 4028 15376
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3700 14816 3752 14822
rect 3620 14764 3700 14770
rect 3620 14758 3752 14764
rect 3344 14634 3372 14758
rect 3620 14742 3740 14758
rect 3344 14618 3464 14634
rect 3240 14612 3292 14618
rect 3344 14612 3476 14618
rect 3344 14606 3424 14612
rect 3240 14554 3292 14560
rect 3424 14554 3476 14560
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2608 12186 2636 12378
rect 1400 12164 1452 12170
rect 1400 12106 1452 12112
rect 2516 12158 2636 12186
rect 2700 12170 2728 13194
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12306 2912 12786
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2688 12164 2740 12170
rect 1412 11762 1440 12106
rect 2516 12102 2544 12158
rect 2688 12106 2740 12112
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 1964 11762 1992 12038
rect 2424 11898 2452 12038
rect 2884 11898 2912 12242
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2976 11558 3004 12106
rect 3068 11830 3096 14350
rect 3240 13932 3292 13938
rect 3344 13920 3372 14486
rect 3620 14414 3648 14742
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3712 14414 3740 14554
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3804 13938 3832 15302
rect 3988 15162 4016 15370
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3988 14414 4016 15098
rect 4172 15026 4200 15422
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14414 4752 15846
rect 4816 15366 4844 16050
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 4816 14618 4844 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5368 15094 5396 15302
rect 5552 15162 5580 16118
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 5000 14414 5028 14758
rect 5092 14618 5304 14634
rect 5080 14612 5304 14618
rect 5132 14606 5304 14612
rect 5080 14554 5132 14560
rect 5276 14550 5304 14606
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 3976 14408 4028 14414
rect 4068 14408 4120 14414
rect 3976 14350 4028 14356
rect 4066 14376 4068 14385
rect 4712 14408 4764 14414
rect 4120 14376 4122 14385
rect 4712 14350 4764 14356
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4066 14311 4122 14320
rect 4816 13938 4844 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 3292 13892 3372 13920
rect 3792 13932 3844 13938
rect 3240 13874 3292 13880
rect 3792 13874 3844 13880
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3160 12170 3188 13806
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 3344 13190 3372 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5000 13326 5028 13670
rect 5276 13530 5304 13942
rect 5368 13938 5396 14418
rect 5552 14414 5580 15098
rect 5644 14822 5672 16662
rect 5828 16250 5856 17614
rect 5920 17066 5948 18142
rect 6288 17746 6316 18566
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6380 17202 6408 19468
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6564 18766 6592 19314
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6472 18358 6500 18634
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 6196 16590 6224 17070
rect 6184 16584 6236 16590
rect 6288 16572 6316 17138
rect 6564 16998 6592 17614
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6656 16726 6684 21014
rect 6748 20874 6776 21422
rect 7024 21298 7052 21490
rect 7116 21418 7144 21966
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 7024 21270 7144 21298
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6840 20058 6868 20742
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6840 19786 6868 19994
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6932 19378 6960 19654
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6368 16584 6420 16590
rect 6288 16544 6368 16572
rect 6184 16526 6236 16532
rect 6368 16526 6420 16532
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 14958 5764 15438
rect 5828 15094 5856 16186
rect 6196 16182 6224 16526
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6380 16114 6408 16526
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5920 15570 5948 15914
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5644 14278 5672 14758
rect 5920 14385 5948 15506
rect 6564 15502 6592 15846
rect 6748 15706 6776 18770
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17882 6960 18226
rect 7024 18222 7052 19110
rect 7116 18222 7144 21270
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7392 20602 7420 20742
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7392 18766 7420 20538
rect 7760 19922 7788 22510
rect 7852 21894 7880 22578
rect 7944 21894 7972 22646
rect 7840 21888 7892 21894
rect 7840 21830 7892 21836
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7472 19236 7524 19242
rect 7472 19178 7524 19184
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6840 17762 6868 17818
rect 6840 17734 7052 17762
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 15700 6788 15706
rect 6656 15660 6736 15688
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6656 15026 6684 15660
rect 6736 15642 6788 15648
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 5906 14376 5962 14385
rect 5816 14340 5868 14346
rect 5906 14311 5962 14320
rect 5816 14282 5868 14288
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4988 13320 5040 13326
rect 5368 13308 5396 13738
rect 5460 13462 5488 14214
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5448 13456 5500 13462
rect 5448 13398 5500 13404
rect 5368 13280 5488 13308
rect 4988 13262 5040 13268
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5460 12850 5488 13280
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12170 3464 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 3068 11150 3096 11766
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10742 3096 11086
rect 3252 11082 3280 12038
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 11354 3464 11766
rect 3620 11626 3648 12310
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3712 11898 3740 12038
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3620 10810 3648 11562
rect 3804 11082 3832 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3896 11558 3924 11766
rect 3988 11762 4016 11834
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 4080 11234 4108 12038
rect 4448 11830 4476 12174
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4632 11558 4660 12786
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 11762 4752 12582
rect 4816 11898 4844 12718
rect 5460 12238 5488 12786
rect 5552 12714 5580 13874
rect 5644 13802 5672 14214
rect 5828 13938 5856 14282
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5828 13734 5856 13874
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5644 12442 5672 13262
rect 5736 12850 5764 13262
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11898 5304 12106
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 4802 11792 4858 11801
rect 4712 11756 4764 11762
rect 4802 11727 4858 11736
rect 5170 11792 5226 11801
rect 5368 11778 5396 12038
rect 5276 11762 5396 11778
rect 5170 11727 5172 11736
rect 4712 11698 4764 11704
rect 4816 11694 4844 11727
rect 5224 11727 5226 11736
rect 5264 11756 5396 11762
rect 5172 11698 5224 11704
rect 5316 11750 5396 11756
rect 5264 11698 5316 11704
rect 4804 11688 4856 11694
rect 4856 11648 4936 11676
rect 4804 11630 4856 11636
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4080 11206 4292 11234
rect 4724 11218 4752 11562
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11354 4844 11494
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4908 11234 4936 11648
rect 4264 11150 4292 11206
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4816 11206 4936 11234
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 3804 10810 3832 11018
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 3068 10062 3096 10678
rect 4172 10674 4200 10950
rect 4356 10742 4384 11018
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1780 8634 1808 9590
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1964 8566 1992 9114
rect 2608 8634 2636 9454
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8974 2820 9318
rect 2976 8974 3004 9386
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7342 1992 8230
rect 2608 7818 2636 8570
rect 2976 8498 3004 8910
rect 3056 8560 3108 8566
rect 3240 8560 3292 8566
rect 3108 8508 3240 8514
rect 3056 8502 3292 8508
rect 2964 8492 3016 8498
rect 3068 8486 3280 8502
rect 2964 8434 3016 8440
rect 2780 8424 2832 8430
rect 2832 8372 3280 8378
rect 2780 8366 3280 8372
rect 2792 8350 3280 8366
rect 3252 8294 3280 8350
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3160 8090 3188 8230
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2332 7410 2360 7686
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 6866 1992 7278
rect 2608 6914 2636 7754
rect 2516 6886 2636 6914
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 5370 1992 6802
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6390 2176 6598
rect 2332 6458 2360 6666
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2516 6118 2544 6886
rect 2792 6458 2820 8026
rect 3344 8022 3372 9318
rect 3436 8838 3464 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3436 7342 3464 8774
rect 3528 7886 3556 9114
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3620 8566 3648 9046
rect 4724 8974 4752 9998
rect 4816 9382 4844 11206
rect 5276 11150 5304 11698
rect 5356 11688 5408 11694
rect 5460 11642 5488 12174
rect 5408 11636 5488 11642
rect 5356 11630 5488 11636
rect 5368 11614 5488 11630
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5368 10962 5396 11614
rect 5644 11558 5672 12242
rect 5736 11898 5764 12786
rect 5828 12102 5856 12854
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5276 10934 5396 10962
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 8968 4764 8974
rect 4526 8936 4582 8945
rect 4908 8922 4936 9386
rect 4712 8910 4764 8916
rect 4816 8906 4936 8922
rect 4526 8871 4582 8880
rect 4620 8900 4672 8906
rect 4540 8566 4568 8871
rect 4620 8842 4672 8848
rect 4816 8900 4948 8906
rect 4816 8894 4896 8900
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 3620 7886 3648 8502
rect 4632 8294 4660 8842
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3528 7750 3556 7822
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3528 7206 3556 7686
rect 3620 7478 3648 7822
rect 3804 7546 3832 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3252 6798 3280 7142
rect 3620 6866 3648 7414
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3896 6798 3924 7822
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 3160 6322 3188 6666
rect 3252 6322 3280 6734
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 6322 3740 6598
rect 4080 6458 4108 7822
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7546 4384 7754
rect 4632 7750 4660 8230
rect 4724 7886 4752 8774
rect 4816 8498 4844 8894
rect 4896 8842 4948 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8566 5304 10934
rect 5552 10742 5580 11290
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5644 10470 5672 11494
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 10810 5764 11018
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5920 9674 5948 14311
rect 6012 13938 6040 14962
rect 6656 14890 6684 14962
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6104 14482 6132 14758
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6564 14414 6592 14758
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6012 13802 6040 13874
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 6196 13462 6224 14350
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6472 14006 6500 14214
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6288 13530 6316 13942
rect 6656 13870 6684 14350
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6748 13716 6776 15302
rect 6656 13688 6776 13716
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6196 12986 6224 13398
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5736 9646 5948 9674
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5460 8974 5488 9114
rect 5736 8974 5764 9646
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 5908 9104 5960 9110
rect 6184 9104 6236 9110
rect 5960 9064 6184 9092
rect 5908 9046 5960 9052
rect 6184 9046 6236 9052
rect 6472 8974 6500 9114
rect 6564 9042 6592 9318
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 5448 8968 5500 8974
rect 5724 8968 5776 8974
rect 5448 8910 5500 8916
rect 5630 8936 5686 8945
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5276 7886 5304 8502
rect 5460 8294 5488 8910
rect 5540 8900 5592 8906
rect 6460 8968 6512 8974
rect 5724 8910 5776 8916
rect 6182 8936 6238 8945
rect 5630 8871 5632 8880
rect 5540 8842 5592 8848
rect 5684 8871 5686 8880
rect 5908 8900 5960 8906
rect 5632 8842 5684 8848
rect 6460 8910 6512 8916
rect 6182 8871 6238 8880
rect 5908 8842 5960 8848
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5552 8022 5580 8842
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8090 5672 8434
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5736 7954 5764 8774
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5828 8090 5856 8570
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5828 7750 5856 7890
rect 5920 7886 5948 8842
rect 6196 8634 6224 8871
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 4632 7546 4660 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 5552 7478 5580 7686
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6798 4660 7346
rect 5828 6798 5856 7686
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 2608 6202 2636 6258
rect 2608 6174 2728 6202
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2516 5914 2544 6054
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1964 4690 1992 5306
rect 2516 5098 2544 5850
rect 2608 5642 2636 6054
rect 2700 5710 2728 6174
rect 3160 5710 3188 6258
rect 3436 6186 3464 6258
rect 4172 6186 4200 6734
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6390 4660 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4436 5908 4488 5914
rect 4632 5896 4660 6326
rect 5276 5914 5304 6326
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5552 5914 5580 6054
rect 4488 5868 4660 5896
rect 5264 5908 5316 5914
rect 4436 5850 4488 5856
rect 5264 5850 5316 5856
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 2608 5098 2636 5578
rect 2700 5234 2728 5646
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5370 3280 5510
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 2240 4622 2268 4966
rect 2700 4842 2728 5170
rect 4448 5030 4476 5850
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4632 5098 4660 5238
rect 5276 5234 5304 5646
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5552 5370 5580 5578
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 5736 5030 5764 6054
rect 5828 5370 5856 6734
rect 6104 6322 6132 7958
rect 6380 7818 6408 8230
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6472 6458 6500 8230
rect 6656 7886 6684 13688
rect 6840 13326 6868 16934
rect 7024 13530 7052 17734
rect 7116 17202 7144 18158
rect 7208 17814 7236 18226
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7300 17678 7328 18294
rect 7392 17746 7420 18362
rect 7484 18086 7512 19178
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7208 17542 7236 17614
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17202 7236 17478
rect 7104 17196 7156 17202
rect 7104 17138 7156 17144
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7392 15502 7420 17682
rect 7576 17542 7604 18566
rect 7760 18222 7788 19858
rect 7852 19446 7880 21830
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7944 19242 7972 21830
rect 8220 21554 8248 21830
rect 8312 21622 8340 23054
rect 8496 22642 8524 23258
rect 8680 22710 8708 23462
rect 10520 23322 10548 23666
rect 10508 23316 10560 23322
rect 10508 23258 10560 23264
rect 10888 23186 10916 23666
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 11072 23050 11100 24550
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11164 23089 11192 23598
rect 11150 23080 11206 23089
rect 8760 23044 8812 23050
rect 8760 22986 8812 22992
rect 11060 23044 11112 23050
rect 11150 23015 11152 23024
rect 11060 22986 11112 22992
rect 11204 23015 11206 23024
rect 11152 22986 11204 22992
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8312 20874 8340 21558
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8312 20534 8340 20810
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8404 20058 8432 20810
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8496 19990 8524 22578
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7852 18290 7880 18838
rect 8128 18426 8156 19178
rect 8220 18465 8248 19382
rect 8206 18456 8262 18465
rect 8116 18420 8168 18426
rect 8206 18391 8262 18400
rect 8116 18362 8168 18368
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7760 17814 7788 18158
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7944 17678 7972 18294
rect 8220 18222 8248 18391
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8312 17746 8340 19926
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8404 18834 8432 19314
rect 8496 19310 8524 19790
rect 8588 19666 8616 22578
rect 8680 22166 8708 22646
rect 8772 22506 8800 22986
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 8760 22500 8812 22506
rect 8760 22442 8812 22448
rect 8668 22160 8720 22166
rect 8668 22102 8720 22108
rect 9048 20874 9076 22918
rect 11072 22574 11100 22986
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 11152 22094 11204 22098
rect 11256 22094 11284 23598
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11348 23186 11376 23462
rect 11440 23254 11468 24142
rect 11716 23322 11744 24142
rect 11808 23866 11836 24686
rect 11900 24138 11928 24754
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11900 23866 11928 24074
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11704 23316 11756 23322
rect 11704 23258 11756 23264
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11612 23248 11664 23254
rect 11612 23190 11664 23196
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11624 22778 11652 23190
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11992 22642 12020 23258
rect 12084 23254 12112 24754
rect 13188 24682 13216 26930
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12164 23724 12216 23730
rect 12164 23666 12216 23672
rect 12176 23322 12204 23666
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 12084 22574 12112 23054
rect 12268 22624 12296 24006
rect 12360 23798 12388 24142
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12360 23118 12388 23734
rect 12452 23322 12480 23802
rect 12544 23730 12572 24278
rect 13188 24138 13216 24618
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13280 24410 13308 24550
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 13372 24070 13400 24686
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12452 22710 12480 23258
rect 12544 23118 12572 23666
rect 13372 23662 13400 24006
rect 13360 23656 13412 23662
rect 13360 23598 13412 23604
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 13004 23118 13032 23462
rect 13096 23186 13124 23462
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13372 23118 13400 23598
rect 13556 23497 13584 23598
rect 13820 23520 13872 23526
rect 13542 23488 13598 23497
rect 13820 23462 13872 23468
rect 13542 23423 13598 23432
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13740 23118 13768 23258
rect 13832 23186 13860 23462
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 12532 23112 12584 23118
rect 12716 23112 12768 23118
rect 12532 23054 12584 23060
rect 12714 23080 12716 23089
rect 12992 23112 13044 23118
rect 12768 23080 12770 23089
rect 12992 23054 13044 23060
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 12714 23015 12770 23024
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22778 13216 22986
rect 13372 22982 13400 23054
rect 13360 22976 13412 22982
rect 13360 22918 13412 22924
rect 13728 22976 13780 22982
rect 13924 22930 13952 24754
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 14016 23322 14044 23666
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14292 23089 14320 24550
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 17592 24200 17644 24206
rect 18144 24200 18196 24206
rect 17644 24160 17724 24188
rect 17592 24142 17644 24148
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16764 24064 16816 24070
rect 16764 24006 16816 24012
rect 14476 23798 14504 24006
rect 14464 23792 14516 23798
rect 14464 23734 14516 23740
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14278 23080 14334 23089
rect 14278 23015 14334 23024
rect 13780 22924 13952 22930
rect 13728 22918 13952 22924
rect 13740 22902 13952 22918
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12268 22596 12388 22624
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 11152 22092 11284 22094
rect 11204 22066 11284 22092
rect 11152 22034 11204 22040
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9140 21690 9168 21966
rect 11164 21894 11192 22034
rect 11440 22030 11468 22510
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8680 19854 8708 20198
rect 8956 19922 8984 20810
rect 9140 20534 9168 21626
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9496 21344 9548 21350
rect 9496 21286 9548 21292
rect 9508 21078 9536 21286
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9600 20942 9628 21422
rect 10152 20942 10180 21830
rect 11256 21146 11284 21966
rect 11716 21962 11744 22374
rect 11900 22030 11928 22374
rect 11888 22024 11940 22030
rect 11808 21984 11888 22012
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21554 11744 21898
rect 11808 21690 11836 21984
rect 11888 21966 11940 21972
rect 11888 21888 11940 21894
rect 11888 21830 11940 21836
rect 11900 21690 11928 21830
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11992 21554 12020 22374
rect 12084 21554 12112 22510
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12268 22166 12296 22442
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12268 21690 12296 22102
rect 12360 22030 12388 22596
rect 13832 22438 13860 22902
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11992 21146 12020 21490
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 9324 20602 9352 20742
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 9128 20528 9180 20534
rect 11532 20505 11560 20742
rect 9128 20470 9180 20476
rect 11518 20496 11574 20505
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9048 19854 9076 20470
rect 11518 20431 11574 20440
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10520 19854 10548 20334
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 8668 19712 8720 19718
rect 8588 19660 8668 19666
rect 8588 19654 8720 19660
rect 8588 19638 8708 19654
rect 8680 19310 8708 19638
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8496 18902 8524 19246
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8404 18630 8432 18770
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18426 8432 18566
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7576 17202 7604 17478
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7668 16998 7696 17478
rect 8496 17134 8524 18022
rect 8588 17338 8616 18226
rect 8680 17610 8708 19246
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8772 17746 8800 18566
rect 8850 18456 8906 18465
rect 8850 18391 8852 18400
rect 8904 18391 8906 18400
rect 8852 18362 8904 18368
rect 8956 17814 8984 18702
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9692 17882 9720 18634
rect 10140 18216 10192 18222
rect 10244 18204 10272 18702
rect 10336 18358 10364 19110
rect 10428 18358 10456 19178
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10324 18352 10376 18358
rect 10324 18294 10376 18300
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10520 18222 10548 18906
rect 10796 18902 10824 19110
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10192 18176 10272 18204
rect 10140 18158 10192 18164
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8956 17202 8984 17750
rect 10060 17678 10088 18022
rect 10244 17678 10272 18176
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 11072 17610 11100 19790
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11440 19378 11468 19722
rect 11532 19378 11560 19790
rect 11900 19786 11928 20742
rect 12084 19854 12112 21490
rect 12360 21468 12388 21966
rect 12176 21440 12388 21468
rect 12176 20942 12204 21440
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 12268 18698 12296 21286
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12452 20534 12480 20878
rect 12544 20602 12572 21966
rect 12820 21690 12848 21966
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12716 21616 12768 21622
rect 12716 21558 12768 21564
rect 12728 21146 12756 21558
rect 12820 21146 12848 21626
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12714 21040 12770 21049
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12636 20534 12664 21014
rect 12714 20975 12716 20984
rect 12768 20975 12770 20984
rect 12716 20946 12768 20952
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12820 20641 12848 20878
rect 12806 20632 12862 20641
rect 12912 20602 12940 21490
rect 13082 21040 13138 21049
rect 12992 21004 13044 21010
rect 13082 20975 13138 20984
rect 12992 20946 13044 20952
rect 12806 20567 12862 20576
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12452 19514 12480 20470
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12452 19394 12480 19450
rect 12360 19366 12480 19394
rect 12360 18834 12388 19366
rect 12544 18970 12572 20198
rect 12912 19854 12940 20334
rect 13004 20262 13032 20946
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 13096 19334 13124 20975
rect 13188 20466 13216 21830
rect 13556 21690 13584 21966
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 13464 21146 13492 21558
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13464 21010 13584 21026
rect 13648 21010 13676 21286
rect 13726 21040 13782 21049
rect 13452 21004 13584 21010
rect 13504 20998 13584 21004
rect 13452 20946 13504 20952
rect 13450 20496 13506 20505
rect 13176 20460 13228 20466
rect 13556 20466 13584 20998
rect 13636 21004 13688 21010
rect 13726 20975 13782 20984
rect 13636 20946 13688 20952
rect 13450 20431 13452 20440
rect 13176 20402 13228 20408
rect 13504 20431 13506 20440
rect 13544 20460 13596 20466
rect 13452 20402 13504 20408
rect 13544 20402 13596 20408
rect 13556 20346 13584 20402
rect 13372 20330 13584 20346
rect 13360 20324 13584 20330
rect 13412 20318 13584 20324
rect 13360 20266 13412 20272
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13096 19306 13216 19334
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 10980 17134 11008 17546
rect 11072 17338 11100 17546
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13938 7512 14214
rect 7668 13938 7696 14962
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6840 12782 6868 13262
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 7300 12646 7328 13738
rect 7484 13530 7512 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 11354 6776 11698
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6748 11082 6776 11290
rect 7208 11082 7236 12242
rect 7300 11354 7328 12582
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7378 11112 7434 11121
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 7196 11076 7248 11082
rect 7378 11047 7380 11056
rect 7196 11018 7248 11024
rect 7432 11047 7434 11056
rect 7380 11018 7432 11024
rect 7104 10736 7156 10742
rect 7208 10724 7236 11018
rect 7484 10810 7512 13262
rect 7760 12918 7788 13874
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 13326 7880 13670
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7852 12986 7880 13262
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7668 11082 7696 11630
rect 7852 11354 7880 11698
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 10810 7696 11018
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7156 10696 7236 10724
rect 7104 10678 7156 10684
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 8838 6776 10542
rect 7944 9110 7972 17070
rect 10980 16046 11008 17070
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 14006 8064 14350
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13530 8064 13806
rect 8128 13802 8156 14554
rect 8588 14414 8616 15438
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8300 14000 8352 14006
rect 8352 13960 8432 13988
rect 8300 13942 8352 13948
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8312 13394 8340 13670
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12850 8064 13126
rect 8128 12986 8156 13262
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 8036 11218 8064 11698
rect 8220 11694 8248 13194
rect 8404 12986 8432 13960
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13190 8524 13806
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8588 12918 8616 14350
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8772 13530 8800 13942
rect 8852 13932 8904 13938
rect 8956 13920 8984 15302
rect 8904 13892 8984 13920
rect 8852 13874 8904 13880
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 12986 8708 13194
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8496 12238 8524 12786
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8312 11354 8340 12174
rect 8496 11898 8524 12174
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 11014 8064 11154
rect 8312 11150 8340 11290
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8208 11144 8260 11150
rect 8206 11112 8208 11121
rect 8300 11144 8352 11150
rect 8260 11112 8262 11121
rect 8300 11086 8352 11092
rect 8206 11047 8262 11056
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8496 10742 8524 11222
rect 8588 11218 8616 12854
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8680 11082 8708 12038
rect 8772 11830 8800 12174
rect 8864 11880 8892 13874
rect 9048 13734 9076 15370
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9140 13938 9168 14962
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8956 12442 8984 12854
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 9048 12306 9076 13670
rect 9140 13394 9168 13874
rect 9232 13734 9260 14962
rect 9600 14618 9628 15370
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15026 10272 15302
rect 10980 15094 11008 15982
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11624 15026 11652 16390
rect 11716 16182 11744 18566
rect 11900 18086 11928 18566
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 12084 17814 12112 18634
rect 12452 18426 12480 18838
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12268 18290 12296 18362
rect 12544 18306 12572 18906
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12360 18278 12572 18306
rect 13004 18290 13032 18566
rect 13096 18426 13124 18702
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13188 18290 13216 19306
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 12360 18222 12388 18278
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12544 18086 12572 18278
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12544 17882 12572 18022
rect 12636 17882 12664 18158
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16794 11836 17138
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 12268 16658 12296 16934
rect 12452 16658 12480 17478
rect 12912 17202 12940 18090
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12912 16998 12940 17138
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12452 16250 12480 16594
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11716 15706 11744 16118
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11808 15026 11836 15846
rect 12084 15706 12112 16050
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12268 15502 12296 15846
rect 12820 15638 12848 16390
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12912 15570 12940 16390
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 15094 12388 15438
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9784 14414 9812 14962
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14482 11376 14758
rect 11624 14618 11652 14962
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11808 14414 11836 14962
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 14414 12020 14486
rect 13004 14482 13032 16458
rect 13176 15496 13228 15502
rect 13096 15444 13176 15450
rect 13096 15438 13228 15444
rect 13096 15422 13216 15438
rect 13096 15026 13124 15422
rect 13280 15162 13308 19246
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13372 17882 13400 18770
rect 13464 18358 13492 20198
rect 13648 19310 13676 20946
rect 13740 20942 13768 20975
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13832 20602 13860 21286
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13648 18766 13676 19246
rect 13832 19242 13860 19654
rect 13924 19514 13952 22646
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14002 20632 14058 20641
rect 14002 20567 14004 20576
rect 14056 20567 14058 20576
rect 14004 20538 14056 20544
rect 14108 20534 14136 21082
rect 14292 21010 14320 23015
rect 14568 22982 14596 23666
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14660 21894 14688 23190
rect 14752 22778 14780 23666
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15580 23118 15608 23462
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15476 22432 15528 22438
rect 15476 22374 15528 22380
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14108 19854 14136 20470
rect 14292 20262 14320 20946
rect 14384 20466 14412 21014
rect 14476 21010 14504 21830
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14844 21146 14872 21490
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15028 20534 15056 20878
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20602 15240 20742
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13542 18456 13598 18465
rect 13542 18391 13544 18400
rect 13596 18391 13598 18400
rect 13544 18362 13596 18368
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13648 18222 13676 18702
rect 13832 18426 13860 18906
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 14016 18290 14044 19110
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 14108 17882 14136 19314
rect 14384 18290 14412 20402
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14476 20058 14504 20334
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14476 19514 14504 19994
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19514 14872 19722
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15212 18834 15240 20198
rect 15304 19310 15332 20266
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14476 18426 14504 18702
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14568 17610 14596 18702
rect 15212 17882 15240 18770
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 16998 14596 17546
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13372 15706 13400 16050
rect 13648 16046 13676 16594
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13648 15570 13676 15982
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15162 13400 15302
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13372 15026 13400 15098
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9324 13938 9352 14214
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9312 13184 9364 13190
rect 9416 13172 9444 13942
rect 9508 13326 9536 13942
rect 9600 13734 9628 14214
rect 11808 13938 11836 14350
rect 11992 14090 12020 14350
rect 11992 14062 12112 14090
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 11796 13932 11848 13938
rect 11848 13892 12020 13920
rect 11796 13874 11848 13880
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9364 13144 9444 13172
rect 9312 13126 9364 13132
rect 9324 12646 9352 13126
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9324 12238 9352 12582
rect 9508 12306 9536 13262
rect 9600 13258 9628 13670
rect 10060 13530 10088 13874
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12306 11008 12718
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 8864 11852 8984 11880
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8864 11354 8892 11698
rect 8956 11558 8984 11852
rect 10980 11762 11008 12242
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 11286 8984 11494
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 10980 10742 11008 11698
rect 11808 11354 11836 11698
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9692 9926 9720 10610
rect 10980 10062 11008 10678
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10130 11284 10610
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6840 8430 6868 8910
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6644 7880 6696 7886
rect 6840 7868 6868 8230
rect 7208 7886 7236 9046
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8634 9076 8774
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 6920 7880 6972 7886
rect 6840 7840 6920 7868
rect 6644 7822 6696 7828
rect 6920 7822 6972 7828
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6564 6458 6592 7822
rect 6656 7546 6684 7822
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 7116 7410 7144 7686
rect 7300 7410 7328 8230
rect 7392 8090 7420 8502
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7546 7420 8026
rect 8036 7750 8064 8366
rect 8772 7750 8800 8570
rect 9324 8498 9352 8910
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9600 8362 9628 9454
rect 9692 8566 9720 9862
rect 9968 9178 9996 9862
rect 10980 9586 11008 9998
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10244 8838 10272 9522
rect 11072 9382 11100 9930
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 10244 8362 10272 8774
rect 10520 8430 10548 8842
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8036 7546 8064 7686
rect 9140 7546 9168 7754
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 10428 7410 10456 7890
rect 10520 7886 10548 8366
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10980 7954 11008 8191
rect 11072 8022 11100 9318
rect 11256 8838 11284 10066
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11256 8430 11284 8774
rect 11348 8634 11376 8774
rect 11532 8634 11560 8910
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11256 7886 11284 8366
rect 11532 8090 11560 8570
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 7852 7002 7880 7346
rect 7944 7274 7972 7346
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6472 6322 6500 6394
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6104 5710 6132 6258
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 5370 6132 5646
rect 6472 5574 6500 6258
rect 6564 5846 6592 6394
rect 7760 6322 7788 6598
rect 7944 6390 7972 7210
rect 8128 6662 8156 7346
rect 8496 7206 8524 7346
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6458 8156 6598
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6564 5386 6592 5782
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6472 5358 6592 5386
rect 6472 5302 6500 5358
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6656 5030 6684 5510
rect 7484 5302 7512 6258
rect 7760 5642 7788 6258
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7944 5302 7972 6326
rect 8312 6118 8340 6326
rect 8496 6322 8524 7142
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8404 6186 8432 6258
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5846 8340 6054
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7944 5098 7972 5238
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 2700 4826 2820 4842
rect 2700 4820 2832 4826
rect 2700 4814 2780 4820
rect 2780 4762 2832 4768
rect 8312 4622 8340 5782
rect 8404 4826 8432 6122
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4690 8524 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8588 5370 8616 5850
rect 8772 5778 8800 6734
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8864 6458 8892 6666
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8956 5914 8984 6258
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8680 5234 8708 5510
rect 8772 5302 8800 5714
rect 9324 5642 9352 6258
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5642 9536 6054
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 10428 2650 10456 7346
rect 10520 6730 10548 7822
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10876 7404 10928 7410
rect 10980 7392 11008 7754
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 10928 7364 11008 7392
rect 10876 7346 10928 7352
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10520 5710 10548 6666
rect 10980 6458 11008 6802
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10968 6316 11020 6322
rect 11072 6304 11100 6870
rect 11348 6798 11376 7210
rect 11440 7002 11468 7686
rect 11532 7410 11560 8026
rect 11624 7546 11652 8434
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 8090 11836 8230
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11716 7410 11744 7890
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11900 7342 11928 13670
rect 11992 7460 12020 13892
rect 12084 13734 12112 14062
rect 12176 14006 12204 14418
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12360 13682 12388 14214
rect 12636 13870 12664 14282
rect 13096 13938 13124 14962
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12440 13728 12492 13734
rect 12360 13676 12440 13682
rect 12360 13670 12492 13676
rect 12360 13654 12480 13670
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 11082 12112 13126
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12360 10810 12388 13654
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 11898 12480 13262
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12452 10674 12480 11018
rect 12636 10674 12664 11086
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 8566 12112 10474
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 9654 12204 10406
rect 12268 10266 12296 10610
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12452 9994 12480 10610
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 12164 9648 12216 9654
rect 12164 9590 12216 9596
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9042 12204 9318
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12452 8838 12480 9930
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 7818 12112 8502
rect 12164 8288 12216 8294
rect 12162 8256 12164 8265
rect 12216 8256 12218 8265
rect 12162 8191 12218 8200
rect 12360 7818 12388 8774
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7834 12480 8230
rect 12544 7954 12572 8774
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12728 8294 12756 8570
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12624 7880 12676 7886
rect 12452 7818 12572 7834
rect 12624 7822 12676 7828
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12348 7812 12400 7818
rect 12452 7812 12584 7818
rect 12452 7806 12532 7812
rect 12348 7754 12400 7760
rect 12532 7754 12584 7760
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 12452 7478 12480 7686
rect 12440 7472 12492 7478
rect 11992 7432 12112 7460
rect 12084 7342 12112 7432
rect 12440 7414 12492 7420
rect 11888 7336 11940 7342
rect 11610 7304 11666 7313
rect 11888 7278 11940 7284
rect 12072 7336 12124 7342
rect 12440 7336 12492 7342
rect 12072 7278 12124 7284
rect 12438 7304 12440 7313
rect 12492 7304 12494 7313
rect 11610 7239 11612 7248
rect 11664 7239 11666 7248
rect 11612 7210 11664 7216
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11900 6730 11928 7278
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 7002 12020 7142
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11020 6276 11100 6304
rect 10968 6258 11020 6264
rect 11348 6254 11376 6598
rect 12084 6390 12112 7278
rect 12438 7239 12494 7248
rect 12636 7002 12664 7822
rect 12728 7410 12756 8230
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5710 10824 6054
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11992 5574 12020 6190
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 11992 2446 12020 5510
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4078 12572 4558
rect 12820 4486 12848 13874
rect 13372 13394 13400 14962
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13556 13326 13584 14214
rect 13648 13870 13676 15370
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14482 13952 14758
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 14016 13530 14044 14962
rect 14752 14074 14780 17274
rect 15212 16658 15240 17818
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15304 15910 15332 16594
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 15570 15332 15846
rect 15396 15570 15424 20402
rect 15488 19310 15516 22374
rect 15580 22030 15608 22510
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15580 19122 15608 21966
rect 15672 21554 15700 23054
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 16040 22642 16068 22918
rect 16224 22778 16252 23598
rect 16500 23186 16528 23734
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16592 23118 16620 24006
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16132 22098 16160 22578
rect 16684 22574 16712 23462
rect 16776 23322 16804 24006
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 22098 16712 22510
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16672 22092 16724 22098
rect 16672 22034 16724 22040
rect 16776 21962 16804 23258
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 22574 17080 22918
rect 17224 22704 17276 22710
rect 17276 22652 17356 22658
rect 17224 22646 17356 22652
rect 17236 22630 17356 22646
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 17052 22030 17080 22510
rect 17328 22166 17356 22630
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 17236 21894 17264 21966
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15672 19922 15700 21490
rect 17328 20942 17356 22102
rect 17604 22030 17632 22510
rect 17696 22506 17724 24160
rect 18144 24142 18196 24148
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17788 23118 17816 23462
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 17880 22438 17908 24006
rect 18156 23798 18184 24142
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 17960 23724 18012 23730
rect 18012 23684 18092 23712
rect 17960 23666 18012 23672
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17972 22710 18000 22918
rect 18064 22778 18092 23684
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 17868 22432 17920 22438
rect 17868 22374 17920 22380
rect 17880 22234 17908 22374
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17972 22094 18000 22646
rect 18340 22642 18368 24074
rect 18708 23712 18736 24142
rect 19156 23724 19208 23730
rect 18708 23684 19012 23712
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 18616 22710 18644 22986
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18708 22642 18736 23462
rect 18984 23118 19012 23684
rect 19156 23666 19208 23672
rect 19168 23322 19196 23666
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18984 22642 19012 23054
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18984 22234 19012 22578
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18052 22094 18104 22098
rect 17972 22092 18104 22094
rect 17972 22066 18052 22092
rect 18052 22034 18104 22040
rect 19076 22030 19104 22918
rect 19168 22642 19196 23122
rect 19156 22636 19208 22642
rect 19260 22624 19288 24210
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23118 19472 24006
rect 19628 23322 19656 24074
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19628 22710 19656 23258
rect 19720 23254 19748 24142
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19616 22704 19668 22710
rect 19616 22646 19668 22652
rect 19340 22636 19392 22642
rect 19260 22596 19340 22624
rect 19156 22578 19208 22584
rect 19340 22578 19392 22584
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 17592 22024 17644 22030
rect 17592 21966 17644 21972
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19076 21010 19104 21966
rect 19168 21350 19196 22374
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19352 22094 19380 22170
rect 19444 22166 19472 22510
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19260 22066 19380 22094
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19310 15700 19858
rect 16684 19854 16712 20742
rect 17420 20602 17448 20946
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15488 19094 15608 19122
rect 15488 18170 15516 19094
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18358 15608 18566
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15672 18272 15700 19246
rect 16684 18970 16712 19314
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 17144 18834 17172 19994
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15752 18284 15804 18290
rect 15672 18244 15752 18272
rect 15752 18226 15804 18232
rect 15488 18142 15608 18170
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15488 17202 15516 17614
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 14822 14872 15302
rect 15200 14952 15252 14958
rect 15396 14906 15424 15506
rect 15200 14894 15252 14900
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 15212 14346 15240 14894
rect 15304 14878 15424 14906
rect 15580 14890 15608 18142
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15948 16794 15976 17478
rect 16040 17202 16068 18566
rect 16868 18086 16896 18702
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16132 17134 16160 17682
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16592 17338 16620 17614
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16868 16658 16896 18022
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 16960 16658 16988 17206
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15568 14884 15620 14890
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15304 14278 15332 14878
rect 15568 14826 15620 14832
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15396 14278 15424 14758
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 11354 12940 12786
rect 13004 11762 13032 13194
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13096 11898 13124 12242
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 13096 11286 13124 11834
rect 13280 11762 13308 12582
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13188 11150 13216 11562
rect 13280 11218 13308 11698
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13176 11144 13228 11150
rect 13372 11098 13400 12174
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 13648 11150 13676 11766
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13176 11086 13228 11092
rect 13188 10810 13216 11086
rect 13280 11070 13400 11098
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9178 12940 9318
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13280 8922 13308 11070
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13740 10062 13768 10542
rect 13360 10056 13412 10062
rect 13728 10056 13780 10062
rect 13360 9998 13412 10004
rect 13648 10016 13728 10044
rect 13188 8894 13308 8922
rect 13188 5234 13216 8894
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8498 13308 8774
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13280 7954 13308 8434
rect 13372 8362 13400 9998
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13464 7954 13492 9862
rect 13648 9178 13676 10016
rect 13728 9998 13780 10004
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 8498 13584 8842
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13648 8430 13676 8910
rect 13740 8430 13768 9318
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8634 13860 8910
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7342 13492 7890
rect 13924 7732 13952 11698
rect 14200 11694 14228 12038
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14200 11354 14228 11494
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14200 10266 14228 11290
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8498 14136 9318
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14200 7886 14228 8502
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 13924 7704 14044 7732
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13832 5846 13860 6734
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13280 4622 13308 4966
rect 13832 4826 13860 5578
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12820 2774 12848 4422
rect 13832 3942 13860 4762
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13740 3534 13768 3878
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13740 3058 13768 3470
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 12636 2746 12848 2774
rect 12636 2514 12664 2746
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13832 2446 13860 3878
rect 13924 2446 13952 6054
rect 14016 5778 14044 7704
rect 14292 7002 14320 13194
rect 14752 12434 14780 14010
rect 15384 14000 15436 14006
rect 15106 13968 15162 13977
rect 15672 13977 15700 14350
rect 15384 13942 15436 13948
rect 15658 13968 15714 13977
rect 15106 13903 15108 13912
rect 15160 13903 15162 13912
rect 15108 13874 15160 13880
rect 15396 13530 15424 13942
rect 15658 13903 15714 13912
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 14660 12406 14780 12434
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11762 14504 12038
rect 14568 11898 14596 12106
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14568 10674 14596 11018
rect 14660 10742 14688 12406
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14752 11762 14780 12174
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14752 11218 14780 11698
rect 14844 11354 14872 12174
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14924 11280 14976 11286
rect 14844 11228 14924 11234
rect 14844 11222 14976 11228
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14844 11206 14964 11222
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14568 10266 14596 10610
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14568 10062 14596 10202
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14660 9518 14688 9862
rect 14752 9586 14780 11154
rect 14844 10674 14872 11206
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10810 14964 10950
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9648 15160 9654
rect 15212 9636 15240 9930
rect 15160 9608 15240 9636
rect 15108 9590 15160 9596
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14568 8498 14596 9454
rect 14752 9042 14780 9522
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14752 8566 14780 8978
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14556 8492 14608 8498
rect 14384 8452 14556 8480
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14108 5914 14136 6258
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5846 14228 6394
rect 14292 6118 14320 6666
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14108 5234 14136 5578
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 5114 14136 5170
rect 14016 5086 14136 5114
rect 14200 5098 14228 5782
rect 14188 5092 14240 5098
rect 14016 4486 14044 5086
rect 14188 5034 14240 5040
rect 14384 4622 14412 8452
rect 14556 8434 14608 8440
rect 15212 8090 15240 9608
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5710 14504 6122
rect 14568 5710 14596 6598
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14476 5370 14504 5646
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14476 4622 14504 5306
rect 14568 4622 14596 5510
rect 14660 5302 14688 6734
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 5846 14780 6190
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14752 5710 14780 5782
rect 15120 5710 15148 6734
rect 15304 5914 15332 13194
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11762 15608 12038
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10810 15424 11018
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15672 10606 15700 11494
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 9994 15700 10542
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9654 15424 9862
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7478 15608 7754
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15396 6458 15424 7346
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6390 15516 6734
rect 15580 6730 15608 7414
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15580 6322 15608 6666
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15382 5808 15438 5817
rect 15580 5778 15608 6258
rect 15382 5743 15438 5752
rect 15568 5772 15620 5778
rect 15396 5710 15424 5743
rect 15568 5714 15620 5720
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4826 14688 5102
rect 14752 4826 14780 5646
rect 15120 5234 15148 5646
rect 15382 5536 15438 5545
rect 15382 5471 15438 5480
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15396 5030 15424 5471
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14752 4622 14780 4762
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14016 2446 14044 4422
rect 14108 4146 14136 4422
rect 14384 4146 14412 4558
rect 14752 4282 14780 4558
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 15396 4146 15424 4966
rect 15488 4826 15516 5170
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15580 4706 15608 5714
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15488 4678 15608 4706
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14384 3466 14412 3878
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 15120 3126 15148 3878
rect 15304 3126 15332 4014
rect 15488 3534 15516 4678
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15580 3194 15608 4082
rect 15672 4010 15700 5646
rect 15764 5234 15792 15030
rect 15856 14074 15884 16390
rect 16960 16114 16988 16594
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 15162 15976 15302
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14346 16712 14758
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16224 13394 16252 14010
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16040 11558 16068 12038
rect 16592 11558 16620 12038
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10606 15976 10950
rect 16488 10804 16540 10810
rect 16488 10746 16540 10752
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 9654 16436 10406
rect 16500 9926 16528 10746
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16500 9518 16528 9862
rect 16488 9512 16540 9518
rect 16408 9460 16488 9466
rect 16408 9454 16540 9460
rect 16408 9438 16528 9454
rect 16580 9444 16632 9450
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 6322 15884 7686
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15948 6458 15976 6598
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16040 6322 16068 6598
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15856 5914 15884 6258
rect 15948 6118 15976 6258
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15856 5370 15884 5578
rect 16132 5574 16160 6938
rect 16408 6338 16436 9438
rect 16580 9386 16632 9392
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 8974 16528 9318
rect 16592 9178 16620 9386
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16684 8498 16712 10678
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16592 7546 16620 7686
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16684 7449 16712 8434
rect 16776 7546 16804 14894
rect 16960 14414 16988 16050
rect 17144 15094 17172 18566
rect 17236 17814 17264 19314
rect 17328 18834 17356 20402
rect 17512 20058 17540 20878
rect 19168 20874 19196 21286
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20466 18736 20742
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 18064 19854 18092 20334
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18064 19310 18092 19790
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17328 17678 17356 18770
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17880 17882 17908 18634
rect 18064 18272 18092 19246
rect 18144 18284 18196 18290
rect 18064 18244 18144 18272
rect 18144 18226 18196 18232
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 18340 17746 18368 19654
rect 19076 19514 19104 19858
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18616 18290 18644 18566
rect 19076 18290 19104 19450
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17604 17270 17632 17546
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 17880 17202 17908 17614
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17880 15910 17908 17138
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15586 17908 15846
rect 17880 15570 18000 15586
rect 17880 15564 18012 15570
rect 17880 15558 17960 15564
rect 17960 15506 18012 15512
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 17144 14550 17172 15030
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17328 14618 17356 14826
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13938 16988 14350
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16868 12306 16896 13874
rect 16960 13394 16988 13874
rect 18248 13530 18276 17478
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18340 16658 18368 17070
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18340 16250 18368 16594
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18340 13410 18368 13738
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 18248 13382 18368 13410
rect 18248 13326 18276 13382
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 12986 17908 13194
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 18248 12782 18276 13262
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17328 11830 17356 12038
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17052 11218 17080 11698
rect 17408 11552 17460 11558
rect 17460 11500 17540 11506
rect 17408 11494 17540 11500
rect 17420 11478 17540 11494
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10674 17172 10950
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16670 7440 16726 7449
rect 16868 7410 16896 8434
rect 17040 7948 17092 7954
rect 17040 7890 17092 7896
rect 16670 7375 16726 7384
rect 16856 7404 16908 7410
rect 16684 6798 16712 7375
rect 16856 7346 16908 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16868 6866 16896 7346
rect 16960 7206 16988 7346
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16856 6724 16908 6730
rect 16960 6712 16988 7142
rect 16908 6684 16988 6712
rect 16856 6666 16908 6672
rect 16408 6310 16528 6338
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15844 5364 15896 5370
rect 16132 5352 16160 5510
rect 15844 5306 15896 5312
rect 16040 5324 16160 5352
rect 16040 5234 16068 5324
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 4146 15884 5102
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4146 16068 4558
rect 16224 4554 16252 6122
rect 16408 5234 16436 6190
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15948 2990 15976 4014
rect 16132 3738 16160 4490
rect 16224 4146 16252 4490
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3754 16436 4082
rect 16500 3942 16528 6310
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16776 5778 16804 6258
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16776 4690 16804 5714
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16408 3738 16528 3754
rect 16120 3732 16172 3738
rect 16408 3732 16540 3738
rect 16408 3726 16488 3732
rect 16120 3674 16172 3680
rect 16488 3674 16540 3680
rect 16132 3126 16160 3674
rect 16592 3126 16620 3946
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16684 3194 16712 3402
rect 16776 3194 16804 4150
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15212 2446 15240 2858
rect 16132 2446 16160 3062
rect 16868 2446 16896 6666
rect 17052 6322 17080 7890
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16960 5846 16988 6258
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 5302 17080 5510
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 3398 16988 4082
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16946 3088 17002 3097
rect 16946 3023 16948 3032
rect 17000 3023 17002 3032
rect 16948 2994 17000 3000
rect 17052 2922 17080 4422
rect 17144 3097 17172 10610
rect 17420 8090 17448 11018
rect 17512 9994 17540 11478
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17420 6118 17448 8026
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5642 17264 5782
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17130 3088 17186 3097
rect 17130 3023 17186 3032
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 17236 2446 17264 5578
rect 17420 4282 17448 5578
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17328 3194 17356 4082
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17420 3058 17448 4218
rect 17512 4146 17540 9930
rect 17604 9518 17632 9998
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17604 8566 17632 9454
rect 17788 9382 17816 12038
rect 18432 11354 18460 17206
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18524 16794 18552 17002
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18524 15638 18552 16730
rect 18708 16590 18736 16934
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 19168 16522 19196 20810
rect 19260 20466 19288 22066
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20534 19472 20742
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19352 19990 19380 20402
rect 19444 20058 19472 20470
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 19718 19288 19790
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19444 19446 19472 19994
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19260 17678 19288 19314
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19352 17882 19380 18362
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19444 17270 19472 18158
rect 19536 17746 19564 22374
rect 19628 22234 19656 22646
rect 19616 22228 19668 22234
rect 19616 22170 19668 22176
rect 19720 21962 19748 23190
rect 20180 23118 20208 24006
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 19812 22438 19840 23054
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19720 20942 19748 21898
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19812 21729 19840 21830
rect 19798 21720 19854 21729
rect 19798 21655 19854 21664
rect 19904 21486 19932 21830
rect 19996 21554 20024 22374
rect 20180 22234 20208 23054
rect 20272 23050 20300 23462
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22692 20300 22986
rect 20352 22704 20404 22710
rect 20272 22664 20352 22692
rect 20352 22646 20404 22652
rect 20364 22506 20392 22646
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 20364 22098 20392 22442
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20548 21672 20576 23122
rect 20640 23050 20668 23666
rect 21008 23186 21036 23666
rect 21100 23322 21128 24074
rect 21192 23662 21220 24550
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 21468 23866 21496 24074
rect 21744 24070 21772 24754
rect 23388 24200 23440 24206
rect 23388 24142 23440 24148
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21456 23860 21508 23866
rect 21456 23802 21508 23808
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21192 23118 21220 23598
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21272 23248 21324 23254
rect 21272 23190 21324 23196
rect 21284 23118 21312 23190
rect 21180 23112 21232 23118
rect 21178 23080 21180 23089
rect 21272 23112 21324 23118
rect 21232 23080 21234 23089
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20812 23044 20864 23050
rect 21272 23054 21324 23060
rect 21178 23015 21234 23024
rect 20812 22986 20864 22992
rect 20626 22944 20682 22953
rect 20626 22879 20682 22888
rect 20640 22030 20668 22879
rect 20824 22778 20852 22986
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20732 22166 20760 22374
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20456 21644 20576 21672
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19996 21146 20024 21354
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20180 20942 20208 21286
rect 20364 20942 20392 21422
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 20168 20936 20220 20942
rect 20352 20936 20404 20942
rect 20168 20878 20220 20884
rect 20350 20904 20352 20913
rect 20404 20904 20406 20913
rect 19720 20466 19748 20878
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19812 20602 19840 20742
rect 19904 20641 19932 20878
rect 19890 20632 19946 20641
rect 19800 20596 19852 20602
rect 19890 20567 19946 20576
rect 19800 20538 19852 20544
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19904 20398 19932 20567
rect 20180 20466 20208 20878
rect 20350 20839 20406 20848
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19800 20324 19852 20330
rect 19800 20266 19852 20272
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19628 18290 19656 18566
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19812 17882 19840 20266
rect 19904 19854 19932 20334
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19904 18329 19932 19790
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 19890 18320 19946 18329
rect 19890 18255 19892 18264
rect 19944 18255 19946 18264
rect 20168 18284 20220 18290
rect 19892 18226 19944 18232
rect 20168 18226 20220 18232
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19800 17876 19852 17882
rect 19800 17818 19852 17824
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17270 19748 17478
rect 19432 17264 19484 17270
rect 19432 17206 19484 17212
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19984 16584 20036 16590
rect 20088 16574 20116 18090
rect 20036 16546 20116 16574
rect 19984 16526 20036 16532
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19720 16114 19748 16458
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 18708 15502 18736 15846
rect 20180 15502 20208 18226
rect 20272 18222 20300 18566
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20272 16794 20300 17138
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20364 16674 20392 20198
rect 20456 18272 20484 21644
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 20330 20576 21490
rect 20732 21486 20760 22102
rect 20824 22030 20852 22578
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 21008 21944 21036 22374
rect 21100 22148 21128 22442
rect 21192 22438 21220 22918
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21180 22160 21232 22166
rect 21100 22120 21180 22148
rect 21180 22102 21232 22108
rect 21008 21916 21128 21944
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20720 21480 20772 21486
rect 20626 21448 20682 21457
rect 20720 21422 20772 21428
rect 20824 21434 20852 21830
rect 20994 21720 21050 21729
rect 20994 21655 21050 21664
rect 21008 21622 21036 21655
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21100 21434 21128 21916
rect 21192 21894 21220 22102
rect 21284 22098 21312 23054
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 21376 22234 21404 22374
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 21554 21220 21830
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21284 21434 21312 21490
rect 20824 21406 20944 21434
rect 20626 21383 20682 21392
rect 20640 21078 20668 21383
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20628 21072 20680 21078
rect 20628 21014 20680 21020
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 20640 20602 20668 20878
rect 20732 20874 20760 21082
rect 20824 20942 20852 21286
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20732 20398 20760 20810
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20824 20058 20852 20878
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20536 18284 20588 18290
rect 20456 18244 20536 18272
rect 20456 18086 20484 18244
rect 20536 18226 20588 18232
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20548 17066 20576 17818
rect 20640 17202 20668 18362
rect 20732 18329 20760 18702
rect 20718 18320 20774 18329
rect 20916 18290 20944 21406
rect 21008 21406 21128 21434
rect 21192 21418 21312 21434
rect 21180 21412 21312 21418
rect 21008 20942 21036 21406
rect 21232 21406 21312 21412
rect 21180 21354 21232 21360
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21008 19990 21036 20878
rect 21100 20398 21128 21286
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 20996 19984 21048 19990
rect 20996 19926 21048 19932
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21008 19514 21036 19790
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 21008 18873 21036 19450
rect 21100 19258 21128 20334
rect 21192 19922 21220 21082
rect 21284 20942 21312 21286
rect 21376 21078 21404 21898
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21284 20330 21312 20878
rect 21376 20777 21404 20878
rect 21362 20768 21418 20777
rect 21362 20703 21418 20712
rect 21362 20632 21418 20641
rect 21362 20567 21364 20576
rect 21416 20567 21418 20576
rect 21364 20538 21416 20544
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21376 19990 21404 20538
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21100 19230 21220 19258
rect 21192 19174 21220 19230
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20994 18864 21050 18873
rect 20994 18799 21050 18808
rect 20718 18255 20720 18264
rect 20772 18255 20774 18264
rect 20904 18284 20956 18290
rect 20720 18226 20772 18232
rect 20904 18226 20956 18232
rect 20916 17746 20944 18226
rect 21008 17882 21036 18799
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20916 17202 20944 17682
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17218 21036 17614
rect 21100 17338 21128 19110
rect 21178 18592 21234 18601
rect 21178 18527 21234 18536
rect 21192 18222 21220 18527
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21192 17610 21220 18158
rect 21284 18086 21312 19654
rect 21376 18630 21404 19790
rect 21468 18766 21496 22374
rect 21560 22234 21588 23258
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22574 21680 23054
rect 21744 23050 21772 24006
rect 23400 23474 23428 24142
rect 23400 23446 23520 23474
rect 22192 23248 22244 23254
rect 22192 23190 22244 23196
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21732 23044 21784 23050
rect 21732 22986 21784 22992
rect 21744 22953 21772 22986
rect 21730 22944 21786 22953
rect 21730 22879 21786 22888
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21548 22002 21600 22008
rect 21548 21944 21600 21950
rect 21560 20874 21588 21944
rect 21652 21486 21680 22510
rect 21732 21548 21784 21554
rect 21836 21536 21864 23054
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22778 21956 22918
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 21928 22094 21956 22170
rect 22100 22094 22152 22098
rect 22204 22094 22232 23190
rect 23492 22642 23520 23446
rect 25228 23112 25280 23118
rect 25228 23054 25280 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25240 22642 25268 23054
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25608 22642 25636 22918
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 23492 22522 23520 22578
rect 23492 22494 23612 22522
rect 21928 22066 22048 22094
rect 22020 21978 22048 22066
rect 22100 22092 22232 22094
rect 22152 22066 22232 22092
rect 22100 22034 22152 22040
rect 22020 21950 22140 21978
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22020 21554 22048 21830
rect 21784 21508 21864 21536
rect 21732 21490 21784 21496
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21836 21418 21864 21508
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21652 20466 21680 21014
rect 21732 20936 21784 20942
rect 21730 20904 21732 20913
rect 21784 20904 21786 20913
rect 21730 20839 21786 20848
rect 21822 20632 21878 20641
rect 21822 20567 21878 20576
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21652 19854 21680 20402
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21652 19446 21680 19790
rect 21836 19718 21864 20567
rect 21928 20466 21956 21490
rect 22008 20800 22060 20806
rect 22006 20768 22008 20777
rect 22060 20768 22062 20777
rect 22006 20703 22062 20712
rect 22006 20632 22062 20641
rect 22006 20567 22062 20576
rect 22020 20482 22048 20567
rect 22112 20482 22140 21950
rect 22204 21690 22232 22066
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22204 20534 22232 21626
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22296 21146 22324 21558
rect 22388 21457 22416 21830
rect 22374 21448 22430 21457
rect 22374 21383 22430 21392
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22284 20868 22336 20874
rect 22284 20810 22336 20816
rect 22020 20466 22140 20482
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 21916 20460 21968 20466
rect 22020 20460 22152 20466
rect 22020 20454 22100 20460
rect 21916 20402 21968 20408
rect 22100 20402 22152 20408
rect 21928 20058 21956 20402
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21640 19440 21692 19446
rect 21640 19382 21692 19388
rect 21928 19378 21956 19994
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21560 18766 21588 19110
rect 21456 18760 21508 18766
rect 21454 18728 21456 18737
rect 21548 18760 21600 18766
rect 21508 18728 21510 18737
rect 21548 18702 21600 18708
rect 21730 18728 21786 18737
rect 21454 18663 21510 18672
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 21284 17610 21312 17818
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20904 17196 20956 17202
rect 21008 17190 21128 17218
rect 21284 17202 21312 17546
rect 21376 17338 21404 18090
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 20904 17138 20956 17144
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20364 16646 20484 16674
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20364 15910 20392 16526
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20272 15434 20300 15846
rect 20364 15638 20392 15846
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 18524 14414 18552 15370
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18616 14618 18644 15302
rect 20456 14958 20484 16646
rect 20548 16590 20576 17002
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20732 15502 20760 17138
rect 21100 17134 21128 17190
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20824 16250 20852 16934
rect 20916 16658 20944 16934
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20904 16516 20956 16522
rect 20904 16458 20956 16464
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20916 16114 20944 16458
rect 21100 16454 21128 17070
rect 21284 16522 21312 17138
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21376 15706 21404 17070
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18524 14074 18552 14350
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18616 14074 18644 14282
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 18984 14074 19012 14214
rect 19812 14074 19840 14214
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19260 12986 19288 13126
rect 19536 12986 19564 13874
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19904 12850 19932 13398
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19076 11694 19104 12718
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11898 19380 12038
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18524 11150 18552 11494
rect 18984 11286 19012 11630
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10062 17908 10406
rect 18432 10062 18460 10542
rect 18984 10266 19012 10610
rect 19076 10606 19104 11630
rect 19260 11354 19288 11698
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 17696 8498 17724 8978
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18708 8566 18736 8842
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 18420 8560 18472 8566
rect 18696 8560 18748 8566
rect 18472 8520 18696 8548
rect 18420 8502 18472 8508
rect 18696 8502 18748 8508
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17696 4554 17724 5782
rect 17788 5778 17816 8298
rect 17880 7886 17908 8502
rect 18420 8424 18472 8430
rect 18800 8378 18828 9998
rect 18984 9586 19012 10202
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9654 19288 9862
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18984 9178 19012 9522
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18984 8430 19012 9114
rect 19352 8974 19380 9386
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19076 8498 19104 8774
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18472 8372 18828 8378
rect 18420 8366 18828 8372
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18432 8350 18828 8366
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 18064 6798 18092 7958
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18616 6798 18644 6870
rect 18708 6798 18736 7414
rect 18800 6798 18828 8350
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19076 7546 19104 7686
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 18880 6860 18932 6866
rect 19076 6848 19104 7482
rect 19260 7410 19288 8026
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19168 7313 19196 7346
rect 19154 7304 19210 7313
rect 19154 7239 19210 7248
rect 19168 7002 19196 7239
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 18880 6802 18932 6808
rect 18984 6820 19104 6848
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17972 4622 18000 6598
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5302 18276 5646
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18064 4826 18092 5170
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17512 4049 17540 4082
rect 17696 4078 17724 4490
rect 18156 4146 18184 5102
rect 18340 4758 18368 5850
rect 18892 4826 18920 6802
rect 18984 6730 19012 6820
rect 19156 6792 19208 6798
rect 19076 6752 19156 6780
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 19076 6254 19104 6752
rect 19156 6734 19208 6740
rect 19352 6390 19380 7142
rect 19444 7002 19472 7346
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19076 5778 19104 6190
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 18892 4622 18920 4762
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18892 4214 18920 4558
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 17684 4072 17736 4078
rect 17498 4040 17554 4049
rect 17684 4014 17736 4020
rect 17498 3975 17554 3984
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3466 17816 3878
rect 18156 3534 18184 4082
rect 18984 3738 19012 4558
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19260 3738 19288 4082
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 18696 3664 18748 3670
rect 18696 3606 18748 3612
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17328 2922 17356 2994
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 17696 2774 17724 3334
rect 18708 3126 18736 3606
rect 19352 3602 19380 5782
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19444 4622 19472 5306
rect 19536 4842 19564 12718
rect 19628 12442 19656 12786
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19720 12238 19748 12786
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19812 10130 19840 12242
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19904 11354 19932 11698
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20088 10810 20116 14010
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20180 12442 20208 13874
rect 20272 13326 20300 14554
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20364 13530 20392 13874
rect 20456 13734 20484 14282
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20456 12850 20484 13670
rect 20732 13410 20760 14214
rect 20824 13530 20852 14486
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20548 13382 20852 13410
rect 20916 13394 20944 13874
rect 20548 13326 20576 13382
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20168 12436 20220 12442
rect 20548 12434 20576 13262
rect 20824 12850 20852 13382
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20720 12640 20772 12646
rect 21008 12594 21036 15302
rect 21468 15026 21496 18226
rect 21560 17678 21588 18702
rect 21730 18663 21786 18672
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21652 18290 21680 18566
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17746 21680 18022
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21652 17202 21680 17682
rect 21744 17678 21772 18663
rect 21824 18624 21876 18630
rect 21928 18612 21956 19314
rect 22020 19174 22048 20266
rect 22204 20058 22232 20334
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 22112 19394 22140 19790
rect 22204 19514 22232 19994
rect 22296 19854 22324 20810
rect 22388 20448 22416 21383
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 20874 22600 21286
rect 22560 20868 22612 20874
rect 22560 20810 22612 20816
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22468 20460 22520 20466
rect 22388 20420 22468 20448
rect 22520 20420 22600 20448
rect 22468 20402 22520 20408
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22112 19366 22232 19394
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 22020 18737 22048 18770
rect 22006 18728 22062 18737
rect 22006 18663 22062 18672
rect 22008 18624 22060 18630
rect 21928 18601 22008 18612
rect 21824 18566 21876 18572
rect 21914 18592 22008 18601
rect 21836 18426 21864 18566
rect 21970 18584 22008 18592
rect 22008 18566 22060 18572
rect 21914 18527 21970 18536
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21836 18290 21864 18362
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21928 17678 21956 18090
rect 22112 18086 22140 19178
rect 22204 18698 22232 19366
rect 22388 18986 22416 19722
rect 22480 19514 22508 19858
rect 22572 19854 22600 20420
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22388 18970 22508 18986
rect 22388 18964 22520 18970
rect 22388 18958 22468 18964
rect 22468 18906 22520 18912
rect 22282 18864 22338 18873
rect 22282 18799 22338 18808
rect 22296 18766 22324 18799
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22192 18692 22244 18698
rect 22192 18634 22244 18640
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21916 17672 21968 17678
rect 21968 17632 22048 17660
rect 21916 17614 21968 17620
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21836 16590 21864 16934
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21928 16522 21956 17478
rect 22020 17202 22048 17632
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21560 16114 21588 16390
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 21744 16046 21772 16390
rect 22020 16114 22048 17138
rect 22112 16726 22140 17274
rect 22204 17066 22232 18634
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22296 17814 22324 18226
rect 22284 17808 22336 17814
rect 22284 17750 22336 17756
rect 22296 17270 22324 17750
rect 22388 17338 22416 18702
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22480 16998 22508 18906
rect 22572 18902 22600 19110
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 22100 16720 22152 16726
rect 22664 16674 22692 20742
rect 22756 18290 22784 22034
rect 23492 21706 23520 22034
rect 23400 21690 23520 21706
rect 23388 21684 23520 21690
rect 23440 21678 23520 21684
rect 23388 21626 23440 21632
rect 23584 21554 23612 22494
rect 24412 22234 24440 22578
rect 24768 22568 24820 22574
rect 25884 22545 25912 23054
rect 24768 22510 24820 22516
rect 25870 22536 25926 22545
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24780 22030 24808 22510
rect 25870 22471 25926 22480
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22940 20942 22968 21422
rect 23216 20942 23244 21490
rect 23676 21418 23704 21898
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23768 21010 23796 21490
rect 23952 21146 23980 21830
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 24044 21146 24072 21490
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 22940 20602 22968 20878
rect 23216 20788 23244 20878
rect 23124 20760 23244 20788
rect 23664 20800 23716 20806
rect 23124 20602 23152 20760
rect 23664 20742 23716 20748
rect 23676 20602 23704 20742
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22744 18284 22796 18290
rect 22744 18226 22796 18232
rect 22756 18154 22784 18226
rect 22744 18148 22796 18154
rect 22744 18090 22796 18096
rect 22100 16662 22152 16668
rect 22480 16646 22692 16674
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21744 15570 21772 15982
rect 21914 15600 21970 15609
rect 21732 15564 21784 15570
rect 21914 15535 21970 15544
rect 21732 15506 21784 15512
rect 21928 15502 21956 15535
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 22020 15162 22048 16050
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22112 15094 22140 16050
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 14074 21128 14350
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 14074 21404 14214
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21638 13968 21694 13977
rect 21638 13903 21640 13912
rect 21692 13903 21694 13912
rect 21640 13874 21692 13880
rect 21744 13802 21772 14758
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20720 12582 20772 12588
rect 20548 12406 20668 12434
rect 20168 12378 20220 12384
rect 20272 12306 20576 12322
rect 20260 12300 20576 12306
rect 20312 12294 20576 12300
rect 20260 12242 20312 12248
rect 20548 12238 20576 12294
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11762 20208 12038
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19984 10532 20036 10538
rect 19984 10474 20036 10480
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19996 9382 20024 10474
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19628 8498 19656 8978
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19996 7834 20024 9318
rect 20088 8498 20116 9590
rect 20180 9586 20208 11698
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20272 10538 20300 11086
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20088 7954 20116 8434
rect 20076 7948 20128 7954
rect 20076 7890 20128 7896
rect 19996 7806 20116 7834
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19812 6322 19840 7346
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19812 6118 19840 6258
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19996 5030 20024 7210
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20088 4842 20116 7806
rect 20272 6254 20300 8570
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 5710 20300 6190
rect 20260 5704 20312 5710
rect 20180 5664 20260 5692
rect 20180 5234 20208 5664
rect 20260 5646 20312 5652
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 19536 4814 19932 4842
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19444 4078 19472 4422
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 3602 19472 4014
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17880 2774 17908 2994
rect 17696 2746 17816 2774
rect 17880 2746 18000 2774
rect 17788 2446 17816 2746
rect 17972 2514 18000 2746
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18340 2446 18368 3062
rect 18800 3058 18828 3402
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 19352 2854 19380 3402
rect 19432 3392 19484 3398
rect 19430 3360 19432 3369
rect 19484 3360 19486 3369
rect 19430 3295 19486 3304
rect 19536 3058 19564 4490
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19628 3194 19656 4218
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19720 3641 19748 3946
rect 19706 3632 19762 3641
rect 19812 3602 19840 4150
rect 19706 3567 19762 3576
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19708 3528 19760 3534
rect 19760 3476 19840 3482
rect 19708 3470 19840 3476
rect 19720 3454 19840 3470
rect 19706 3224 19762 3233
rect 19616 3188 19668 3194
rect 19812 3194 19840 3454
rect 19904 3194 19932 4814
rect 19996 4814 20116 4842
rect 19706 3159 19762 3168
rect 19800 3188 19852 3194
rect 19616 3130 19668 3136
rect 19720 3058 19748 3159
rect 19800 3130 19852 3136
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19996 3074 20024 4814
rect 20180 4282 20208 5170
rect 20272 4622 20300 5170
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20168 4276 20220 4282
rect 20220 4236 20300 4264
rect 20168 4218 20220 4224
rect 20166 4176 20222 4185
rect 20076 4140 20128 4146
rect 20166 4111 20222 4120
rect 20076 4082 20128 4088
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19904 3046 20024 3074
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 18616 2650 18644 2790
rect 19536 2774 19564 2994
rect 19444 2746 19564 2774
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18616 2446 18644 2586
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 10336 800 10364 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 800 11652 2246
rect 12268 800 12296 2382
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 12912 800 12940 2246
rect 13556 800 13584 2246
rect 14200 800 14228 2246
rect 14844 800 14872 2246
rect 15488 800 15516 2246
rect 16132 800 16160 2246
rect 16776 800 16804 2246
rect 17420 800 17448 2246
rect 18064 800 18092 2246
rect 18708 800 18736 2518
rect 19444 2514 19472 2746
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19720 2446 19748 2994
rect 19904 2854 19932 3046
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 20088 2378 20116 4082
rect 20180 3534 20208 4111
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20272 3398 20300 4236
rect 20364 3398 20392 12174
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11150 20484 12038
rect 20548 11558 20576 12174
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20548 11218 20576 11494
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8974 20484 9318
rect 20548 9042 20576 11154
rect 20640 11014 20668 12406
rect 20732 12374 20760 12582
rect 20824 12566 21036 12594
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9518 20668 9998
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20732 9058 20760 11562
rect 20824 9382 20852 12566
rect 21100 12434 21128 13466
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 12986 21220 13194
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21284 12986 21312 13126
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21468 12850 21496 13738
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21560 13530 21588 13670
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21560 13326 21588 13466
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21836 13258 21864 14282
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21928 13530 21956 13874
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 12866 21864 13194
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 21652 12850 21864 12866
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21640 12844 21864 12850
rect 21692 12838 21864 12844
rect 21640 12786 21692 12792
rect 21008 12406 21128 12434
rect 21192 12434 21220 12786
rect 21192 12406 21312 12434
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20916 10130 20944 11766
rect 21008 11014 21036 12406
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20640 9030 20760 9058
rect 20916 9042 20944 10066
rect 21008 10062 21036 10406
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20904 9036 20956 9042
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20456 7478 20484 8910
rect 20640 8022 20668 9030
rect 20904 8978 20956 8984
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20732 8634 20760 8910
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20916 8566 20944 8978
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20904 8560 20956 8566
rect 20824 8520 20904 8548
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20628 8016 20680 8022
rect 20628 7958 20680 7964
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 6186 20576 7346
rect 20628 7200 20680 7206
rect 20732 7154 20760 8230
rect 20824 7886 20852 8520
rect 20904 8502 20956 8508
rect 21008 8362 21036 8570
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20680 7148 20760 7154
rect 20628 7142 20760 7148
rect 20640 7126 20760 7142
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20548 5846 20576 6122
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20456 4146 20484 5170
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20548 4214 20576 5034
rect 20536 4208 20588 4214
rect 20534 4176 20536 4185
rect 20588 4176 20590 4185
rect 20444 4140 20496 4146
rect 20590 4134 20668 4162
rect 20534 4111 20590 4120
rect 20444 4082 20496 4088
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20166 3224 20222 3233
rect 20166 3159 20222 3168
rect 20180 2990 20208 3159
rect 20272 3058 20300 3334
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20168 2984 20220 2990
rect 20168 2926 20220 2932
rect 20364 2582 20392 3130
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 20456 2446 20484 3946
rect 20548 3641 20576 4014
rect 20534 3632 20590 3641
rect 20534 3567 20590 3576
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20548 2854 20576 3470
rect 20640 3126 20668 4134
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20640 2961 20668 3062
rect 20626 2952 20682 2961
rect 20626 2887 20682 2896
rect 20536 2848 20588 2854
rect 20536 2790 20588 2796
rect 20732 2446 20760 6598
rect 20824 6202 20852 7346
rect 20916 7324 20944 8026
rect 20996 7812 21048 7818
rect 20996 7754 21048 7760
rect 21008 7546 21036 7754
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 20996 7336 21048 7342
rect 20916 7296 20996 7324
rect 20996 7278 21048 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6798 20944 7142
rect 21008 6798 21036 7278
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20996 6792 21048 6798
rect 20996 6734 21048 6740
rect 20824 6174 21036 6202
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20824 5302 20852 5578
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 20916 5114 20944 6054
rect 21008 5370 21036 6174
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20824 5086 20944 5114
rect 20824 2774 20852 5086
rect 21008 4826 21036 5306
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20902 3360 20958 3369
rect 20902 3295 20958 3304
rect 20916 3058 20944 3295
rect 21100 3194 21128 12174
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21192 3942 21220 11086
rect 21284 9926 21312 12406
rect 21468 12374 21496 12786
rect 21456 12368 21508 12374
rect 21362 12336 21418 12345
rect 21456 12310 21508 12316
rect 21362 12271 21418 12280
rect 21376 12238 21404 12271
rect 21836 12238 21864 12838
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21364 12232 21416 12238
rect 21824 12232 21876 12238
rect 21364 12174 21416 12180
rect 21638 12200 21694 12209
rect 21376 11898 21404 12174
rect 21824 12174 21876 12180
rect 21638 12135 21694 12144
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21376 11218 21404 11834
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21468 10248 21496 11086
rect 21560 10810 21588 11086
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21548 10260 21600 10266
rect 21468 10220 21548 10248
rect 21548 10202 21600 10208
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 8498 21588 8774
rect 21364 8492 21416 8498
rect 21284 8452 21364 8480
rect 21284 7750 21312 8452
rect 21364 8434 21416 8440
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21284 6798 21312 7686
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21468 6866 21496 7346
rect 21560 7002 21588 8434
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21652 6914 21680 12135
rect 21836 11626 21864 12174
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21928 11354 21956 11698
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21836 10452 21864 11018
rect 21916 10600 21968 10606
rect 22020 10588 22048 12718
rect 22112 12102 22140 13126
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 11150 22140 11494
rect 22204 11286 22232 14554
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 21968 10560 22048 10588
rect 21916 10542 21968 10548
rect 21836 10424 21956 10452
rect 21928 9586 21956 10424
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21836 7478 21864 7754
rect 21824 7472 21876 7478
rect 21822 7440 21824 7449
rect 21876 7440 21878 7449
rect 21822 7375 21878 7384
rect 21928 7324 21956 9522
rect 22020 9518 22048 10560
rect 22296 10198 22324 10746
rect 22388 10674 22416 11086
rect 22376 10668 22428 10674
rect 22376 10610 22428 10616
rect 22284 10192 22336 10198
rect 22284 10134 22336 10140
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 22020 7546 22048 9454
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22112 8498 22140 9046
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21836 7296 21956 7324
rect 21652 6886 21772 6914
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21468 6746 21496 6802
rect 21284 6322 21312 6734
rect 21468 6718 21680 6746
rect 21744 6730 21772 6886
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21284 5574 21312 6258
rect 21376 5642 21404 6598
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21272 5568 21324 5574
rect 21468 5545 21496 6258
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5642 21588 6054
rect 21548 5636 21600 5642
rect 21548 5578 21600 5584
rect 21272 5510 21324 5516
rect 21454 5536 21510 5545
rect 21454 5471 21510 5480
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21284 5234 21312 5306
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21468 4826 21496 5170
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21560 4554 21588 5578
rect 21652 4622 21680 6718
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 6322 21772 6666
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21744 5914 21772 6122
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21744 4826 21772 5170
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21560 4282 21588 4490
rect 21744 4486 21772 4762
rect 21836 4758 21864 7296
rect 22112 6730 22140 7686
rect 22204 7274 22232 8570
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 22112 5574 22140 5850
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 21824 4752 21876 4758
rect 21824 4694 21876 4700
rect 21732 4480 21784 4486
rect 21732 4422 21784 4428
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21008 2854 21036 3062
rect 21192 3058 21220 3334
rect 21376 3058 21404 4082
rect 21468 3233 21496 4150
rect 21560 3534 21588 4218
rect 21744 4146 21772 4422
rect 22112 4282 22140 5306
rect 22204 5302 22232 5646
rect 22192 5296 22244 5302
rect 22192 5238 22244 5244
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22112 4146 22140 4218
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22204 3602 22232 5238
rect 22296 4078 22324 10134
rect 22388 9722 22416 10610
rect 22480 9994 22508 16646
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22572 12209 22600 16050
rect 22664 15978 22692 16050
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22664 15638 22692 15914
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22664 14890 22692 15438
rect 22652 14884 22704 14890
rect 22652 14826 22704 14832
rect 22756 13977 22784 15506
rect 22848 14618 22876 20334
rect 22940 18698 22968 20538
rect 23124 20466 23152 20538
rect 23112 20460 23164 20466
rect 23112 20402 23164 20408
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23124 20262 23152 20402
rect 23112 20256 23164 20262
rect 23112 20198 23164 20204
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22940 16164 22968 18634
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23032 16590 23060 17070
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23020 16176 23072 16182
rect 22940 16136 23020 16164
rect 23020 16118 23072 16124
rect 23124 15978 23152 20198
rect 23308 19990 23336 20402
rect 23296 19984 23348 19990
rect 23296 19926 23348 19932
rect 23584 19718 23612 20402
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23768 19378 23796 20946
rect 25240 20942 25268 21286
rect 25424 21185 25452 21830
rect 25410 21176 25466 21185
rect 25410 21111 25466 21120
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24688 20602 24716 20810
rect 25608 20602 25636 21966
rect 25792 21865 25820 22374
rect 25964 21888 26016 21894
rect 25778 21856 25834 21865
rect 25964 21830 26016 21836
rect 25778 21791 25834 21800
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25792 20466 25820 20742
rect 25976 20505 26004 21830
rect 25962 20496 26018 20505
rect 25780 20460 25832 20466
rect 25962 20431 26018 20440
rect 25780 20402 25832 20408
rect 23940 19848 23992 19854
rect 25320 19848 25372 19854
rect 23940 19790 23992 19796
rect 24122 19816 24178 19825
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23216 18426 23244 18702
rect 23204 18420 23256 18426
rect 23204 18362 23256 18368
rect 23584 17882 23612 18770
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 23308 16998 23336 17138
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 16114 23612 16934
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 23216 14278 23244 16050
rect 23676 15502 23704 18702
rect 23768 18290 23796 19314
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 17678 23796 18226
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23768 17202 23796 17614
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23860 16538 23888 19654
rect 23952 19514 23980 19790
rect 25320 19790 25372 19796
rect 24122 19751 24178 19760
rect 24136 19718 24164 19751
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24412 19446 24440 19654
rect 24400 19440 24452 19446
rect 24400 19382 24452 19388
rect 24504 18970 24532 19654
rect 25332 19514 25360 19790
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24044 17202 24072 17478
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23860 16510 23980 16538
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23848 16448 23900 16454
rect 23848 16390 23900 16396
rect 23768 16250 23796 16390
rect 23860 16250 23888 16390
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23308 15162 23336 15370
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23400 14414 23428 15370
rect 23768 15094 23796 15642
rect 23756 15088 23808 15094
rect 23756 15030 23808 15036
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23400 14074 23428 14350
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23756 14000 23808 14006
rect 22742 13968 22798 13977
rect 23756 13942 23808 13948
rect 22742 13903 22798 13912
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22940 13258 22968 13670
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23216 13258 23244 13398
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12918 22784 13126
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 23216 12434 23244 13194
rect 23216 12406 23336 12434
rect 22652 12232 22704 12238
rect 22558 12200 22614 12209
rect 22652 12174 22704 12180
rect 22558 12135 22614 12144
rect 22664 10810 22692 12174
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22940 11354 22968 12106
rect 23204 12096 23256 12102
rect 23204 12038 23256 12044
rect 23216 11558 23244 12038
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22940 11082 22968 11290
rect 23216 11218 23244 11494
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22388 8974 22416 9658
rect 22836 9104 22888 9110
rect 22836 9046 22888 9052
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22388 7750 22416 8434
rect 22848 8430 22876 9046
rect 22940 8906 22968 11018
rect 23308 10742 23336 12406
rect 23400 12238 23428 13262
rect 23664 13252 23716 13258
rect 23768 13240 23796 13942
rect 23716 13212 23796 13240
rect 23664 13194 23716 13200
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23492 12374 23520 12854
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23584 12442 23612 12786
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11218 23428 12174
rect 23676 11830 23704 12786
rect 23768 12782 23796 13212
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23860 12306 23888 16050
rect 23952 13326 23980 16510
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 24044 13938 24072 14214
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13462 24164 13874
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23940 13184 23992 13190
rect 23940 13126 23992 13132
rect 23952 12850 23980 13126
rect 24044 12850 24072 13262
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24136 12986 24164 13194
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24136 12434 24164 12922
rect 23952 12406 24164 12434
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23664 11620 23716 11626
rect 23664 11562 23716 11568
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23308 9738 23336 10678
rect 23400 10674 23428 11154
rect 23584 10674 23612 11222
rect 23676 11218 23704 11562
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23676 10810 23704 11154
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23308 9710 23428 9738
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23308 9178 23336 9522
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23400 9042 23428 9710
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 22836 8424 22888 8430
rect 22836 8366 22888 8372
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22480 6866 22508 7278
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 22664 6254 22692 7278
rect 22940 6798 22968 8842
rect 23400 8634 23428 8978
rect 23492 8974 23520 9862
rect 23676 9738 23704 10746
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23768 10538 23796 10610
rect 23860 10538 23888 11630
rect 23952 11150 23980 12406
rect 24124 11756 24176 11762
rect 24124 11698 24176 11704
rect 24136 11150 24164 11698
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24228 10674 24256 18634
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24320 17746 24348 18566
rect 24412 18358 24440 18566
rect 24400 18352 24452 18358
rect 24400 18294 24452 18300
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24492 17536 24544 17542
rect 24492 17478 24544 17484
rect 24504 15978 24532 17478
rect 24492 15972 24544 15978
rect 24492 15914 24544 15920
rect 24596 15910 24624 18566
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24780 15978 24808 17070
rect 24768 15972 24820 15978
rect 24768 15914 24820 15920
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24308 15360 24360 15366
rect 24308 15302 24360 15308
rect 24320 15162 24348 15302
rect 24308 15156 24360 15162
rect 24308 15098 24360 15104
rect 24872 14822 24900 19382
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25410 19136 25466 19145
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25148 18426 25176 18702
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25332 18290 25360 19110
rect 25410 19071 25466 19080
rect 25424 18426 25452 19071
rect 25516 18766 25544 19314
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25792 18465 25820 19450
rect 25778 18456 25834 18465
rect 25412 18420 25464 18426
rect 25778 18391 25834 18400
rect 25412 18362 25464 18368
rect 25320 18284 25372 18290
rect 25320 18226 25372 18232
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25148 17338 25176 17614
rect 25608 17338 25636 18226
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25792 17785 25820 18022
rect 25778 17776 25834 17785
rect 25778 17711 25834 17720
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25596 17332 25648 17338
rect 25596 17274 25648 17280
rect 25778 17096 25834 17105
rect 25778 17031 25780 17040
rect 25832 17031 25834 17040
rect 25780 17002 25832 17008
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 26054 16416 26110 16425
rect 25516 16114 25544 16390
rect 26054 16351 26110 16360
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24964 15026 24992 15506
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25240 15162 25268 15438
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25228 15156 25280 15162
rect 25228 15098 25280 15104
rect 25424 15065 25452 15302
rect 25410 15056 25466 15065
rect 24952 15020 25004 15026
rect 25410 14991 25466 15000
rect 24952 14962 25004 14968
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24320 14074 24348 14282
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24412 13977 24440 14350
rect 25700 14278 25728 16050
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25792 15745 25820 15846
rect 25778 15736 25834 15745
rect 26068 15706 26096 16351
rect 25778 15671 25834 15680
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25778 14376 25834 14385
rect 25778 14311 25834 14320
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 24492 14000 24544 14006
rect 24398 13968 24454 13977
rect 24492 13942 24544 13948
rect 24398 13903 24454 13912
rect 24412 13326 24440 13903
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23584 9710 23704 9738
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 22928 6792 22980 6798
rect 22928 6734 22980 6740
rect 23032 6730 23060 8570
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23388 8492 23440 8498
rect 23584 8480 23612 9710
rect 23664 9580 23716 9586
rect 23768 9568 23796 10474
rect 23860 9586 23888 10474
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23716 9540 23796 9568
rect 23848 9580 23900 9586
rect 23664 9522 23716 9528
rect 23848 9522 23900 9528
rect 23860 8498 23888 9522
rect 23440 8452 23612 8480
rect 23756 8492 23808 8498
rect 23388 8434 23440 8440
rect 23124 7886 23152 8434
rect 23492 8362 23520 8452
rect 23756 8434 23808 8440
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23768 8378 23796 8434
rect 23952 8378 23980 9930
rect 24044 9674 24072 9998
rect 24044 9646 24256 9674
rect 23480 8356 23532 8362
rect 23768 8350 24164 8378
rect 23480 8298 23532 8304
rect 23492 7886 23520 8298
rect 23940 7948 23992 7954
rect 23940 7890 23992 7896
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 23124 6474 23152 7822
rect 23296 7472 23348 7478
rect 23296 7414 23348 7420
rect 23308 7313 23336 7414
rect 23492 7410 23520 7822
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23768 7324 23796 7822
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7478 23888 7686
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23952 7410 23980 7890
rect 24032 7812 24084 7818
rect 24032 7754 24084 7760
rect 24044 7410 24072 7754
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23294 7304 23350 7313
rect 23768 7296 23888 7324
rect 23294 7239 23350 7248
rect 23480 7268 23532 7274
rect 23032 6446 23152 6474
rect 23032 6322 23060 6446
rect 23308 6322 23336 7239
rect 23480 7210 23532 7216
rect 23492 6866 23520 7210
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23756 6316 23808 6322
rect 23860 6304 23888 7296
rect 23808 6276 23888 6304
rect 23756 6258 23808 6264
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22572 5953 22600 6190
rect 22558 5944 22614 5953
rect 22558 5879 22614 5888
rect 22664 5710 22692 6190
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 23032 5234 23060 6258
rect 23124 5914 23152 6258
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23032 4622 23060 5170
rect 23216 5166 23244 6258
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 23296 5568 23348 5574
rect 23480 5568 23532 5574
rect 23348 5516 23428 5522
rect 23296 5510 23428 5516
rect 23480 5510 23532 5516
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23308 5494 23428 5510
rect 23296 5296 23348 5302
rect 23296 5238 23348 5244
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23216 4690 23244 4966
rect 23308 4690 23336 5238
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23112 4480 23164 4486
rect 23032 4440 23112 4468
rect 23032 4282 23060 4440
rect 23112 4422 23164 4428
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21454 3224 21510 3233
rect 21454 3159 21510 3168
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21100 2961 21128 2994
rect 21086 2952 21142 2961
rect 21086 2887 21142 2896
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 20824 2746 20944 2774
rect 20916 2514 20944 2746
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 21100 2446 21128 2790
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 21192 2310 21220 2994
rect 21560 2854 21588 3470
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 3194 21864 3402
rect 22204 3194 22232 3538
rect 22480 3534 22508 3878
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22098 3088 22154 3097
rect 22480 3058 22508 3130
rect 22098 3023 22100 3032
rect 22152 3023 22154 3032
rect 22284 3052 22336 3058
rect 22100 2994 22152 3000
rect 22284 2994 22336 3000
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 19444 1170 19472 2246
rect 19352 1142 19472 1170
rect 19352 800 19380 1142
rect 19996 800 20024 2246
rect 20640 800 20668 2246
rect 21284 800 21312 2586
rect 22296 2582 22324 2994
rect 22572 2990 22600 4218
rect 23032 4146 23060 4218
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22848 3398 22876 4082
rect 23124 4026 23152 4218
rect 23032 3998 23152 4026
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22940 3126 22968 3878
rect 23032 3398 23060 3998
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23124 3738 23152 3878
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 22928 3120 22980 3126
rect 22928 3062 22980 3068
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22284 2576 22336 2582
rect 22284 2518 22336 2524
rect 23032 2446 23060 3334
rect 23124 3126 23152 3674
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23216 2446 23244 4626
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23308 4146 23336 4490
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23308 3448 23336 4082
rect 23400 3670 23428 5494
rect 23492 5234 23520 5510
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23676 5098 23704 5510
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23768 4622 23796 5782
rect 23860 5234 23888 6276
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23952 5642 23980 5850
rect 24044 5642 24072 6054
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 24032 5636 24084 5642
rect 24032 5578 24084 5584
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23860 4622 23888 5034
rect 24136 4622 24164 8350
rect 24228 7002 24256 9646
rect 24320 7546 24348 12242
rect 24412 9994 24440 12310
rect 24504 12306 24532 13942
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25056 12442 25084 12786
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25148 12442 25176 12582
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24780 12220 24808 12378
rect 25240 12345 25268 13874
rect 25424 13705 25452 14010
rect 25700 14006 25728 14214
rect 25792 14074 25820 14311
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25410 13696 25466 13705
rect 25410 13631 25466 13640
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25608 12850 25636 13126
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25226 12336 25282 12345
rect 25226 12271 25282 12280
rect 24860 12232 24912 12238
rect 24780 12192 24860 12220
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24596 11082 24624 11766
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24688 10810 24716 12174
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24780 10130 24808 12192
rect 24860 12174 24912 12180
rect 25424 12170 25452 12582
rect 25700 12238 25728 13942
rect 25778 13016 25834 13025
rect 25778 12951 25780 12960
rect 25832 12951 25834 12960
rect 25780 12922 25832 12928
rect 25778 12336 25834 12345
rect 25778 12271 25834 12280
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25608 11762 25636 12038
rect 25792 11898 25820 12271
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25778 11656 25834 11665
rect 25596 11620 25648 11626
rect 25778 11591 25834 11600
rect 25596 11562 25648 11568
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 11150 25360 11494
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24872 10470 24900 11018
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24872 10062 24900 10406
rect 25608 10062 25636 11562
rect 25792 11354 25820 11591
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25778 10976 25834 10985
rect 25778 10911 25834 10920
rect 25792 10810 25820 10911
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25778 10296 25834 10305
rect 25778 10231 25780 10240
rect 25832 10231 25834 10240
rect 25780 10202 25832 10208
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25136 10056 25188 10062
rect 25596 10056 25648 10062
rect 25188 10004 25268 10010
rect 25136 9998 25268 10004
rect 25596 9998 25648 10004
rect 24400 9988 24452 9994
rect 25148 9982 25268 9998
rect 24400 9930 24452 9936
rect 24412 9110 24440 9930
rect 25240 9382 25268 9982
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25424 9625 25452 9862
rect 25410 9616 25466 9625
rect 25410 9551 25466 9560
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 25240 9042 25268 9318
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24504 7886 24532 8774
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24216 6996 24268 7002
rect 24216 6938 24268 6944
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 24596 6798 24624 6938
rect 24688 6934 24716 7346
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24688 6798 24716 6870
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24412 6458 24440 6598
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24596 6304 24624 6734
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24676 6316 24728 6322
rect 24596 6276 24676 6304
rect 24596 5710 24624 6276
rect 24676 6258 24728 6264
rect 24780 6254 24808 6666
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24780 5953 24808 6190
rect 24766 5944 24822 5953
rect 24766 5879 24822 5888
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24780 5642 24808 5879
rect 24872 5710 24900 8298
rect 25056 7546 25084 8842
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6186 24992 6734
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25148 5817 25176 6054
rect 25134 5808 25190 5817
rect 25134 5743 25190 5752
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 23756 4616 23808 4622
rect 23756 4558 23808 4564
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24768 4480 24820 4486
rect 24688 4440 24768 4468
rect 23572 4208 23624 4214
rect 23572 4150 23624 4156
rect 23478 4040 23534 4049
rect 23478 3975 23534 3984
rect 23388 3664 23440 3670
rect 23388 3606 23440 3612
rect 23492 3602 23520 3975
rect 23584 3738 23612 4150
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23846 3632 23902 3641
rect 23480 3596 23532 3602
rect 23846 3567 23902 3576
rect 23480 3538 23532 3544
rect 23860 3466 23888 3567
rect 24688 3534 24716 4440
rect 24768 4422 24820 4428
rect 24872 4146 24900 4490
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24780 3738 24808 4082
rect 24768 3732 24820 3738
rect 24768 3674 24820 3680
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 23480 3460 23532 3466
rect 23308 3420 23480 3448
rect 23308 3194 23336 3420
rect 23480 3402 23532 3408
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23860 3194 23888 3402
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23860 2446 23888 3130
rect 24136 3126 24164 3470
rect 24504 3194 24532 3470
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 25240 3058 25268 8978
rect 25596 8968 25648 8974
rect 25596 8910 25648 8916
rect 25778 8936 25834 8945
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25332 8498 25360 8842
rect 25608 8498 25636 8910
rect 25778 8871 25834 8880
rect 25792 8838 25820 8871
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 26146 8256 26202 8265
rect 26146 8191 26202 8200
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25410 6896 25466 6905
rect 25410 6831 25466 6840
rect 25424 6662 25452 6831
rect 25608 6798 25636 7482
rect 25700 7410 25728 7686
rect 25778 7576 25834 7585
rect 26160 7546 26188 8191
rect 25778 7511 25834 7520
rect 26148 7540 26200 7546
rect 25688 7404 25740 7410
rect 25688 7346 25740 7352
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25412 6656 25464 6662
rect 25412 6598 25464 6604
rect 25608 6390 25636 6734
rect 25792 6662 25820 7511
rect 26148 7482 26200 7488
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25778 6216 25834 6225
rect 25320 6180 25372 6186
rect 25778 6151 25834 6160
rect 25320 6122 25372 6128
rect 25332 5914 25360 6122
rect 25596 6112 25648 6118
rect 25596 6054 25648 6060
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25332 5370 25360 5850
rect 25608 5710 25636 6054
rect 25792 5914 25820 6151
rect 25780 5908 25832 5914
rect 25780 5850 25832 5856
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25504 5636 25556 5642
rect 25504 5578 25556 5584
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25516 4826 25544 5578
rect 25778 5536 25834 5545
rect 25778 5471 25834 5480
rect 25792 5370 25820 5471
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25778 4856 25834 4865
rect 25504 4820 25556 4826
rect 25778 4791 25834 4800
rect 25504 4762 25556 4768
rect 25410 4176 25466 4185
rect 25516 4146 25544 4762
rect 25410 4111 25466 4120
rect 25504 4140 25556 4146
rect 25424 4010 25452 4111
rect 25504 4082 25556 4088
rect 25792 4010 25820 4791
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 25780 4004 25832 4010
rect 25780 3946 25832 3952
rect 25778 3496 25834 3505
rect 25778 3431 25834 3440
rect 25792 3398 25820 3431
rect 25780 3392 25832 3398
rect 25780 3334 25832 3340
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 24872 2446 24900 2994
rect 25780 2848 25832 2854
rect 25778 2816 25780 2825
rect 25832 2816 25834 2825
rect 25778 2751 25834 2760
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 21928 800 21956 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 22572 800 22600 2246
rect 23216 800 23244 2246
rect 23860 800 23888 2246
rect 24504 800 24532 2246
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
<< via2 >>
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 110 25608 166 25664
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 846 21256 902 21312
rect 846 18536 902 18592
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4526 22072 4582 22128
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5078 22072 5134 22128
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 846 15816 902 15872
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4802 19216 4858 19272
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 1490 15000 1546 15056
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4066 14356 4068 14376
rect 4068 14356 4120 14376
rect 4120 14356 4122 14376
rect 4066 14320 4122 14356
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 5906 14320 5962 14376
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4802 11736 4858 11792
rect 5170 11756 5226 11792
rect 5170 11736 5172 11756
rect 5172 11736 5224 11756
rect 5224 11736 5226 11756
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4526 8880 4582 8936
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5630 8900 5686 8936
rect 5630 8880 5632 8900
rect 5632 8880 5684 8900
rect 5684 8880 5686 8900
rect 6182 8880 6238 8936
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 11150 23044 11206 23080
rect 11150 23024 11152 23044
rect 11152 23024 11204 23044
rect 11204 23024 11206 23044
rect 8206 18400 8262 18456
rect 13542 23432 13598 23488
rect 12714 23060 12716 23080
rect 12716 23060 12768 23080
rect 12768 23060 12770 23080
rect 12714 23024 12770 23060
rect 14278 23024 14334 23080
rect 11518 20440 11574 20496
rect 8850 18420 8906 18456
rect 8850 18400 8852 18420
rect 8852 18400 8904 18420
rect 8904 18400 8906 18420
rect 12714 21004 12770 21040
rect 12714 20984 12716 21004
rect 12716 20984 12768 21004
rect 12768 20984 12770 21004
rect 12806 20576 12862 20632
rect 13082 20984 13138 21040
rect 13450 20460 13506 20496
rect 13726 20984 13782 21040
rect 13450 20440 13452 20460
rect 13452 20440 13504 20460
rect 13504 20440 13506 20460
rect 7378 11076 7434 11112
rect 7378 11056 7380 11076
rect 7380 11056 7432 11076
rect 7432 11056 7434 11076
rect 8206 11092 8208 11112
rect 8208 11092 8260 11112
rect 8260 11092 8262 11112
rect 8206 11056 8262 11092
rect 14002 20596 14058 20632
rect 14002 20576 14004 20596
rect 14004 20576 14056 20596
rect 14056 20576 14058 20596
rect 13542 18420 13598 18456
rect 13542 18400 13544 18420
rect 13544 18400 13596 18420
rect 13596 18400 13598 18420
rect 10966 8200 11022 8256
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 12162 8236 12164 8256
rect 12164 8236 12216 8256
rect 12216 8236 12218 8256
rect 12162 8200 12218 8236
rect 11610 7268 11666 7304
rect 12438 7284 12440 7304
rect 12440 7284 12492 7304
rect 12492 7284 12494 7304
rect 11610 7248 11612 7268
rect 11612 7248 11664 7268
rect 11664 7248 11666 7268
rect 12438 7248 12494 7284
rect 15106 13932 15162 13968
rect 15106 13912 15108 13932
rect 15108 13912 15160 13932
rect 15160 13912 15162 13932
rect 15658 13912 15714 13968
rect 15382 5752 15438 5808
rect 15382 5480 15438 5536
rect 16670 7384 16726 7440
rect 16946 3052 17002 3088
rect 16946 3032 16948 3052
rect 16948 3032 17000 3052
rect 17000 3032 17002 3052
rect 17130 3032 17186 3088
rect 19798 21664 19854 21720
rect 21178 23060 21180 23080
rect 21180 23060 21232 23080
rect 21232 23060 21234 23080
rect 21178 23024 21234 23060
rect 20626 22888 20682 22944
rect 20350 20884 20352 20904
rect 20352 20884 20404 20904
rect 20404 20884 20406 20904
rect 19890 20576 19946 20632
rect 20350 20848 20406 20884
rect 19890 18284 19946 18320
rect 19890 18264 19892 18284
rect 19892 18264 19944 18284
rect 19944 18264 19946 18284
rect 20626 21392 20682 21448
rect 20994 21664 21050 21720
rect 20718 18284 20774 18320
rect 21362 20712 21418 20768
rect 21362 20596 21418 20632
rect 21362 20576 21364 20596
rect 21364 20576 21416 20596
rect 21416 20576 21418 20596
rect 20994 18808 21050 18864
rect 20718 18264 20720 18284
rect 20720 18264 20772 18284
rect 20772 18264 20774 18284
rect 21178 18536 21234 18592
rect 21730 22888 21786 22944
rect 21730 20884 21732 20904
rect 21732 20884 21784 20904
rect 21784 20884 21786 20904
rect 21730 20848 21786 20884
rect 21822 20576 21878 20632
rect 22006 20748 22008 20768
rect 22008 20748 22060 20768
rect 22060 20748 22062 20768
rect 22006 20712 22062 20748
rect 22006 20576 22062 20632
rect 22374 21392 22430 21448
rect 21454 18708 21456 18728
rect 21456 18708 21508 18728
rect 21508 18708 21510 18728
rect 21454 18672 21510 18708
rect 19154 7248 19210 7304
rect 17498 3984 17554 4040
rect 21730 18672 21786 18728
rect 22006 18672 22062 18728
rect 21914 18536 21970 18592
rect 22282 18808 22338 18864
rect 25870 22480 25926 22536
rect 21914 15544 21970 15600
rect 21638 13932 21694 13968
rect 21638 13912 21640 13932
rect 21640 13912 21692 13932
rect 21692 13912 21694 13932
rect 19430 3340 19432 3360
rect 19432 3340 19484 3360
rect 19484 3340 19486 3360
rect 19430 3304 19486 3340
rect 19706 3576 19762 3632
rect 19706 3168 19762 3224
rect 20166 4120 20222 4176
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 20534 4156 20536 4176
rect 20536 4156 20588 4176
rect 20588 4156 20590 4176
rect 20534 4120 20590 4156
rect 20166 3168 20222 3224
rect 20534 3576 20590 3632
rect 20626 2896 20682 2952
rect 20902 3304 20958 3360
rect 21362 12280 21418 12336
rect 21638 12144 21694 12200
rect 21822 7420 21824 7440
rect 21824 7420 21876 7440
rect 21876 7420 21878 7440
rect 21822 7384 21878 7420
rect 21454 5480 21510 5536
rect 25410 21120 25466 21176
rect 25778 21800 25834 21856
rect 25962 20440 26018 20496
rect 24122 19760 24178 19816
rect 22742 13912 22798 13968
rect 22558 12144 22614 12200
rect 25410 19080 25466 19136
rect 25778 18400 25834 18456
rect 25778 17720 25834 17776
rect 25778 17060 25834 17096
rect 25778 17040 25780 17060
rect 25780 17040 25832 17060
rect 25832 17040 25834 17060
rect 26054 16360 26110 16416
rect 25410 15000 25466 15056
rect 25778 15680 25834 15736
rect 25778 14320 25834 14376
rect 24398 13912 24454 13968
rect 23294 7248 23350 7304
rect 22558 5888 22614 5944
rect 21454 3168 21510 3224
rect 21086 2896 21142 2952
rect 22098 3052 22154 3088
rect 22098 3032 22100 3052
rect 22100 3032 22152 3052
rect 22152 3032 22154 3052
rect 25410 13640 25466 13696
rect 25226 12280 25282 12336
rect 25778 12980 25834 13016
rect 25778 12960 25780 12980
rect 25780 12960 25832 12980
rect 25832 12960 25834 12980
rect 25778 12280 25834 12336
rect 25778 11600 25834 11656
rect 25778 10920 25834 10976
rect 25778 10260 25834 10296
rect 25778 10240 25780 10260
rect 25780 10240 25832 10260
rect 25832 10240 25834 10260
rect 25410 9560 25466 9616
rect 24766 5888 24822 5944
rect 25134 5752 25190 5808
rect 23478 3984 23534 4040
rect 23846 3576 23902 3632
rect 25778 8880 25834 8936
rect 26146 8200 26202 8256
rect 25410 6840 25466 6896
rect 25778 7520 25834 7576
rect 25778 6160 25834 6216
rect 25778 5480 25834 5536
rect 25778 4800 25834 4856
rect 25410 4120 25466 4176
rect 25778 3440 25834 3496
rect 25778 2796 25780 2816
rect 25780 2796 25832 2816
rect 25832 2796 25834 2816
rect 25778 2760 25834 2796
<< metal3 >>
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 0 25938 800 25968
rect 0 25878 1042 25938
rect 0 25848 800 25878
rect 105 25666 171 25669
rect 982 25666 1042 25878
rect 105 25664 1042 25666
rect 105 25608 110 25664
rect 166 25608 1042 25664
rect 105 25606 1042 25608
rect 105 25603 171 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 13537 23492 13603 23493
rect 13486 23490 13492 23492
rect 13446 23430 13492 23490
rect 13556 23488 13603 23492
rect 13598 23432 13603 23488
rect 13486 23428 13492 23430
rect 13556 23428 13603 23432
rect 13537 23427 13603 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 11145 23082 11211 23085
rect 12709 23082 12775 23085
rect 14273 23082 14339 23085
rect 11145 23080 14339 23082
rect 11145 23024 11150 23080
rect 11206 23024 12714 23080
rect 12770 23024 14278 23080
rect 14334 23024 14339 23080
rect 11145 23022 14339 23024
rect 11145 23019 11211 23022
rect 12709 23019 12775 23022
rect 14273 23019 14339 23022
rect 21173 23084 21239 23085
rect 21173 23080 21220 23084
rect 21284 23082 21290 23084
rect 21173 23024 21178 23080
rect 21173 23020 21220 23024
rect 21284 23022 21330 23082
rect 21284 23020 21290 23022
rect 21173 23019 21239 23020
rect 20621 22946 20687 22949
rect 21725 22946 21791 22949
rect 20621 22944 21791 22946
rect 20621 22888 20626 22944
rect 20682 22888 21730 22944
rect 21786 22888 21791 22944
rect 20621 22886 21791 22888
rect 20621 22883 20687 22886
rect 21725 22883 21791 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 25865 22538 25931 22541
rect 26532 22538 27332 22568
rect 25865 22536 27332 22538
rect 25865 22480 25870 22536
rect 25926 22480 27332 22536
rect 25865 22478 27332 22480
rect 25865 22475 25931 22478
rect 26532 22448 27332 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 4521 22130 4587 22133
rect 5073 22130 5139 22133
rect 4521 22128 5139 22130
rect 4521 22072 4526 22128
rect 4582 22072 5078 22128
rect 5134 22072 5139 22128
rect 4521 22070 5139 22072
rect 4521 22067 4587 22070
rect 5073 22067 5139 22070
rect 25773 21858 25839 21861
rect 26532 21858 27332 21888
rect 25773 21856 27332 21858
rect 25773 21800 25778 21856
rect 25834 21800 27332 21856
rect 25773 21798 27332 21800
rect 25773 21795 25839 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 26532 21768 27332 21798
rect 4870 21727 5186 21728
rect 19793 21722 19859 21725
rect 20989 21722 21055 21725
rect 19793 21720 21055 21722
rect 19793 21664 19798 21720
rect 19854 21664 20994 21720
rect 21050 21664 21055 21720
rect 19793 21662 21055 21664
rect 19793 21659 19859 21662
rect 20989 21659 21055 21662
rect 20621 21450 20687 21453
rect 22369 21450 22435 21453
rect 20621 21448 22435 21450
rect 20621 21392 20626 21448
rect 20682 21392 22374 21448
rect 22430 21392 22435 21448
rect 20621 21390 22435 21392
rect 20621 21387 20687 21390
rect 22369 21387 22435 21390
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 25405 21178 25471 21181
rect 26532 21178 27332 21208
rect 25405 21176 27332 21178
rect 25405 21120 25410 21176
rect 25466 21120 27332 21176
rect 25405 21118 27332 21120
rect 0 21088 800 21118
rect 25405 21115 25471 21118
rect 26532 21088 27332 21118
rect 12709 21042 12775 21045
rect 13077 21042 13143 21045
rect 13721 21042 13787 21045
rect 12709 21040 13787 21042
rect 12709 20984 12714 21040
rect 12770 20984 13082 21040
rect 13138 20984 13726 21040
rect 13782 20984 13787 21040
rect 12709 20982 13787 20984
rect 12709 20979 12775 20982
rect 13077 20979 13143 20982
rect 13721 20979 13787 20982
rect 20345 20906 20411 20909
rect 21725 20906 21791 20909
rect 20345 20904 21791 20906
rect 20345 20848 20350 20904
rect 20406 20848 21730 20904
rect 21786 20848 21791 20904
rect 20345 20846 21791 20848
rect 20345 20843 20411 20846
rect 21725 20843 21791 20846
rect 21357 20770 21423 20773
rect 22001 20772 22067 20773
rect 21950 20770 21956 20772
rect 21357 20768 21834 20770
rect 21357 20712 21362 20768
rect 21418 20712 21834 20768
rect 21357 20710 21834 20712
rect 21910 20710 21956 20770
rect 22020 20768 22067 20772
rect 22062 20712 22067 20768
rect 21357 20707 21423 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 21774 20637 21834 20710
rect 21950 20708 21956 20710
rect 22020 20708 22067 20712
rect 22001 20707 22067 20708
rect 12801 20634 12867 20637
rect 13997 20634 14063 20637
rect 12801 20632 14063 20634
rect 12801 20576 12806 20632
rect 12862 20576 14002 20632
rect 14058 20576 14063 20632
rect 12801 20574 14063 20576
rect 12801 20571 12867 20574
rect 13997 20571 14063 20574
rect 19885 20634 19951 20637
rect 21214 20634 21220 20636
rect 19885 20632 21220 20634
rect 19885 20576 19890 20632
rect 19946 20576 21220 20632
rect 19885 20574 21220 20576
rect 19885 20571 19951 20574
rect 21214 20572 21220 20574
rect 21284 20634 21290 20636
rect 21357 20634 21423 20637
rect 21774 20634 21883 20637
rect 22001 20634 22067 20637
rect 21284 20632 21423 20634
rect 21284 20576 21362 20632
rect 21418 20576 21423 20632
rect 21284 20574 21423 20576
rect 21726 20632 22067 20634
rect 21726 20576 21822 20632
rect 21878 20576 22006 20632
rect 22062 20576 22067 20632
rect 21726 20574 22067 20576
rect 21284 20572 21290 20574
rect 21357 20571 21423 20574
rect 21817 20571 21883 20574
rect 22001 20571 22067 20574
rect 11513 20498 11579 20501
rect 13445 20498 13511 20501
rect 11513 20496 13511 20498
rect 11513 20440 11518 20496
rect 11574 20440 13450 20496
rect 13506 20440 13511 20496
rect 11513 20438 13511 20440
rect 11513 20435 11579 20438
rect 13445 20435 13511 20438
rect 25957 20498 26023 20501
rect 26532 20498 27332 20528
rect 25957 20496 27332 20498
rect 25957 20440 25962 20496
rect 26018 20440 27332 20496
rect 25957 20438 27332 20440
rect 25957 20435 26023 20438
rect 26532 20408 27332 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 24117 19818 24183 19821
rect 26532 19818 27332 19848
rect 24117 19816 27332 19818
rect 24117 19760 24122 19816
rect 24178 19760 27332 19816
rect 24117 19758 27332 19760
rect 24117 19755 24183 19758
rect 26532 19728 27332 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4654 19212 4660 19276
rect 4724 19274 4730 19276
rect 4797 19274 4863 19277
rect 4724 19272 4863 19274
rect 4724 19216 4802 19272
rect 4858 19216 4863 19272
rect 4724 19214 4863 19216
rect 4724 19212 4730 19214
rect 4797 19211 4863 19214
rect 25405 19138 25471 19141
rect 26532 19138 27332 19168
rect 25405 19136 27332 19138
rect 25405 19080 25410 19136
rect 25466 19080 27332 19136
rect 25405 19078 27332 19080
rect 25405 19075 25471 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 26532 19048 27332 19078
rect 4210 19007 4526 19008
rect 20989 18866 21055 18869
rect 22277 18866 22343 18869
rect 20989 18864 22343 18866
rect 20989 18808 20994 18864
rect 21050 18808 22282 18864
rect 22338 18808 22343 18864
rect 20989 18806 22343 18808
rect 20989 18803 21055 18806
rect 22277 18803 22343 18806
rect 21449 18730 21515 18733
rect 21725 18730 21791 18733
rect 22001 18730 22067 18733
rect 21449 18728 22067 18730
rect 21449 18672 21454 18728
rect 21510 18672 21730 18728
rect 21786 18672 22006 18728
rect 22062 18672 22067 18728
rect 21449 18670 22067 18672
rect 21449 18667 21515 18670
rect 21725 18667 21791 18670
rect 22001 18667 22067 18670
rect 841 18594 907 18597
rect 798 18592 907 18594
rect 798 18536 846 18592
rect 902 18536 907 18592
rect 798 18531 907 18536
rect 21173 18594 21239 18597
rect 21909 18594 21975 18597
rect 21173 18592 21975 18594
rect 21173 18536 21178 18592
rect 21234 18536 21914 18592
rect 21970 18536 21975 18592
rect 21173 18534 21975 18536
rect 21173 18531 21239 18534
rect 21909 18531 21975 18534
rect 798 18488 858 18531
rect 0 18398 858 18488
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 8201 18458 8267 18461
rect 8845 18458 8911 18461
rect 13537 18460 13603 18461
rect 8201 18456 8911 18458
rect 8201 18400 8206 18456
rect 8262 18400 8850 18456
rect 8906 18400 8911 18456
rect 8201 18398 8911 18400
rect 0 18368 800 18398
rect 8201 18395 8267 18398
rect 8845 18395 8911 18398
rect 13486 18396 13492 18460
rect 13556 18458 13603 18460
rect 25773 18458 25839 18461
rect 26532 18458 27332 18488
rect 13556 18456 13648 18458
rect 13598 18400 13648 18456
rect 13556 18398 13648 18400
rect 25773 18456 27332 18458
rect 25773 18400 25778 18456
rect 25834 18400 27332 18456
rect 25773 18398 27332 18400
rect 13556 18396 13603 18398
rect 13537 18395 13603 18396
rect 25773 18395 25839 18398
rect 26532 18368 27332 18398
rect 19885 18322 19951 18325
rect 20713 18322 20779 18325
rect 19885 18320 20779 18322
rect 19885 18264 19890 18320
rect 19946 18264 20718 18320
rect 20774 18264 20779 18320
rect 19885 18262 20779 18264
rect 19885 18259 19951 18262
rect 20713 18259 20779 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 25773 17778 25839 17781
rect 26532 17778 27332 17808
rect 25773 17776 27332 17778
rect 25773 17720 25778 17776
rect 25834 17720 27332 17776
rect 25773 17718 27332 17720
rect 25773 17715 25839 17718
rect 26532 17688 27332 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 25773 17098 25839 17101
rect 26532 17098 27332 17128
rect 25773 17096 27332 17098
rect 25773 17040 25778 17096
rect 25834 17040 27332 17096
rect 25773 17038 27332 17040
rect 25773 17035 25839 17038
rect 26532 17008 27332 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 26049 16418 26115 16421
rect 26532 16418 27332 16448
rect 26049 16416 27332 16418
rect 26049 16360 26054 16416
rect 26110 16360 27332 16416
rect 26049 16358 27332 16360
rect 26049 16355 26115 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 26532 16328 27332 16358
rect 4870 16287 5186 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 25773 15738 25839 15741
rect 26532 15738 27332 15768
rect 25773 15736 27332 15738
rect 25773 15680 25778 15736
rect 25834 15680 27332 15736
rect 25773 15678 27332 15680
rect 0 15648 800 15678
rect 25773 15675 25839 15678
rect 26532 15648 27332 15678
rect 21909 15604 21975 15605
rect 21909 15602 21956 15604
rect 21864 15600 21956 15602
rect 21864 15544 21914 15600
rect 21864 15542 21956 15544
rect 21909 15540 21956 15542
rect 22020 15540 22026 15604
rect 21909 15539 21975 15540
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 25405 15058 25471 15061
rect 26532 15058 27332 15088
rect 25405 15056 27332 15058
rect 25405 15000 25410 15056
rect 25466 15000 27332 15056
rect 25405 14998 27332 15000
rect 25405 14995 25471 14998
rect 26532 14968 27332 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4061 14378 4127 14381
rect 5901 14378 5967 14381
rect 4061 14376 5967 14378
rect 4061 14320 4066 14376
rect 4122 14320 5906 14376
rect 5962 14320 5967 14376
rect 4061 14318 5967 14320
rect 4061 14315 4127 14318
rect 5901 14315 5967 14318
rect 25773 14378 25839 14381
rect 26532 14378 27332 14408
rect 25773 14376 27332 14378
rect 25773 14320 25778 14376
rect 25834 14320 27332 14376
rect 25773 14318 27332 14320
rect 25773 14315 25839 14318
rect 26532 14288 27332 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 15101 13970 15167 13973
rect 15653 13970 15719 13973
rect 15101 13968 15719 13970
rect 15101 13912 15106 13968
rect 15162 13912 15658 13968
rect 15714 13912 15719 13968
rect 15101 13910 15719 13912
rect 15101 13907 15167 13910
rect 15653 13907 15719 13910
rect 21633 13970 21699 13973
rect 22737 13970 22803 13973
rect 24393 13970 24459 13973
rect 21633 13968 24459 13970
rect 21633 13912 21638 13968
rect 21694 13912 22742 13968
rect 22798 13912 24398 13968
rect 24454 13912 24459 13968
rect 21633 13910 24459 13912
rect 21633 13907 21699 13910
rect 22737 13907 22803 13910
rect 24393 13907 24459 13910
rect 25405 13698 25471 13701
rect 26532 13698 27332 13728
rect 25405 13696 27332 13698
rect 25405 13640 25410 13696
rect 25466 13640 27332 13696
rect 25405 13638 27332 13640
rect 25405 13635 25471 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 26532 13608 27332 13638
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 25773 13018 25839 13021
rect 26532 13018 27332 13048
rect 25773 13016 27332 13018
rect 25773 12960 25778 13016
rect 25834 12960 27332 13016
rect 25773 12958 27332 12960
rect 25773 12955 25839 12958
rect 26532 12928 27332 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 21357 12338 21423 12341
rect 25221 12338 25287 12341
rect 21357 12336 25287 12338
rect 21357 12280 21362 12336
rect 21418 12280 25226 12336
rect 25282 12280 25287 12336
rect 21357 12278 25287 12280
rect 21357 12275 21423 12278
rect 25221 12275 25287 12278
rect 25773 12338 25839 12341
rect 26532 12338 27332 12368
rect 25773 12336 27332 12338
rect 25773 12280 25778 12336
rect 25834 12280 27332 12336
rect 25773 12278 27332 12280
rect 25773 12275 25839 12278
rect 26532 12248 27332 12278
rect 21633 12202 21699 12205
rect 22553 12202 22619 12205
rect 21633 12200 22619 12202
rect 21633 12144 21638 12200
rect 21694 12144 22558 12200
rect 22614 12144 22619 12200
rect 21633 12142 22619 12144
rect 21633 12139 21699 12142
rect 22553 12139 22619 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4654 11732 4660 11796
rect 4724 11794 4730 11796
rect 4797 11794 4863 11797
rect 5165 11794 5231 11797
rect 4724 11792 5231 11794
rect 4724 11736 4802 11792
rect 4858 11736 5170 11792
rect 5226 11736 5231 11792
rect 4724 11734 5231 11736
rect 4724 11732 4730 11734
rect 4797 11731 4863 11734
rect 5165 11731 5231 11734
rect 25773 11658 25839 11661
rect 26532 11658 27332 11688
rect 25773 11656 27332 11658
rect 25773 11600 25778 11656
rect 25834 11600 27332 11656
rect 25773 11598 27332 11600
rect 25773 11595 25839 11598
rect 26532 11568 27332 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 7373 11114 7439 11117
rect 8201 11114 8267 11117
rect 7373 11112 8267 11114
rect 7373 11056 7378 11112
rect 7434 11056 8206 11112
rect 8262 11056 8267 11112
rect 7373 11054 8267 11056
rect 7373 11051 7439 11054
rect 8201 11051 8267 11054
rect 25773 10978 25839 10981
rect 26532 10978 27332 11008
rect 25773 10976 27332 10978
rect 25773 10920 25778 10976
rect 25834 10920 27332 10976
rect 25773 10918 27332 10920
rect 25773 10915 25839 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 26532 10888 27332 10918
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 25773 10298 25839 10301
rect 26532 10298 27332 10328
rect 25773 10296 27332 10298
rect 25773 10240 25778 10296
rect 25834 10240 27332 10296
rect 25773 10238 27332 10240
rect 25773 10235 25839 10238
rect 26532 10208 27332 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 25405 9618 25471 9621
rect 26532 9618 27332 9648
rect 25405 9616 27332 9618
rect 25405 9560 25410 9616
rect 25466 9560 27332 9616
rect 25405 9558 27332 9560
rect 25405 9555 25471 9558
rect 26532 9528 27332 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4521 8938 4587 8941
rect 5625 8938 5691 8941
rect 6177 8938 6243 8941
rect 4521 8936 6243 8938
rect 4521 8880 4526 8936
rect 4582 8880 5630 8936
rect 5686 8880 6182 8936
rect 6238 8880 6243 8936
rect 4521 8878 6243 8880
rect 4521 8875 4587 8878
rect 5625 8875 5691 8878
rect 6177 8875 6243 8878
rect 25773 8938 25839 8941
rect 26532 8938 27332 8968
rect 25773 8936 27332 8938
rect 25773 8880 25778 8936
rect 25834 8880 27332 8936
rect 25773 8878 27332 8880
rect 25773 8875 25839 8878
rect 26532 8848 27332 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 10961 8258 11027 8261
rect 12157 8258 12223 8261
rect 10961 8256 12223 8258
rect 10961 8200 10966 8256
rect 11022 8200 12162 8256
rect 12218 8200 12223 8256
rect 10961 8198 12223 8200
rect 10961 8195 11027 8198
rect 12157 8195 12223 8198
rect 26141 8258 26207 8261
rect 26532 8258 27332 8288
rect 26141 8256 27332 8258
rect 26141 8200 26146 8256
rect 26202 8200 27332 8256
rect 26141 8198 27332 8200
rect 26141 8195 26207 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 26532 8168 27332 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 25773 7578 25839 7581
rect 26532 7578 27332 7608
rect 25773 7576 27332 7578
rect 25773 7520 25778 7576
rect 25834 7520 27332 7576
rect 25773 7518 27332 7520
rect 25773 7515 25839 7518
rect 26532 7488 27332 7518
rect 16665 7442 16731 7445
rect 21817 7442 21883 7445
rect 16665 7440 21883 7442
rect 16665 7384 16670 7440
rect 16726 7384 21822 7440
rect 21878 7384 21883 7440
rect 16665 7382 21883 7384
rect 16665 7379 16731 7382
rect 21817 7379 21883 7382
rect 11605 7306 11671 7309
rect 12433 7306 12499 7309
rect 11605 7304 12499 7306
rect 11605 7248 11610 7304
rect 11666 7248 12438 7304
rect 12494 7248 12499 7304
rect 11605 7246 12499 7248
rect 11605 7243 11671 7246
rect 12433 7243 12499 7246
rect 19149 7306 19215 7309
rect 23289 7306 23355 7309
rect 19149 7304 23355 7306
rect 19149 7248 19154 7304
rect 19210 7248 23294 7304
rect 23350 7248 23355 7304
rect 19149 7246 23355 7248
rect 19149 7243 19215 7246
rect 23289 7243 23355 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 25405 6898 25471 6901
rect 26532 6898 27332 6928
rect 25405 6896 27332 6898
rect 25405 6840 25410 6896
rect 25466 6840 27332 6896
rect 25405 6838 27332 6840
rect 25405 6835 25471 6838
rect 26532 6808 27332 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 25773 6218 25839 6221
rect 26532 6218 27332 6248
rect 25773 6216 27332 6218
rect 25773 6160 25778 6216
rect 25834 6160 27332 6216
rect 25773 6158 27332 6160
rect 25773 6155 25839 6158
rect 26532 6128 27332 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 22553 5946 22619 5949
rect 24761 5946 24827 5949
rect 22553 5944 24827 5946
rect 22553 5888 22558 5944
rect 22614 5888 24766 5944
rect 24822 5888 24827 5944
rect 22553 5886 24827 5888
rect 22553 5883 22619 5886
rect 24761 5883 24827 5886
rect 15377 5810 15443 5813
rect 25129 5810 25195 5813
rect 15377 5808 25195 5810
rect 15377 5752 15382 5808
rect 15438 5752 25134 5808
rect 25190 5752 25195 5808
rect 15377 5750 25195 5752
rect 15377 5747 15443 5750
rect 25129 5747 25195 5750
rect 15377 5538 15443 5541
rect 21449 5538 21515 5541
rect 15377 5536 21515 5538
rect 15377 5480 15382 5536
rect 15438 5480 21454 5536
rect 21510 5480 21515 5536
rect 15377 5478 21515 5480
rect 15377 5475 15443 5478
rect 21449 5475 21515 5478
rect 25773 5538 25839 5541
rect 26532 5538 27332 5568
rect 25773 5536 27332 5538
rect 25773 5480 25778 5536
rect 25834 5480 27332 5536
rect 25773 5478 27332 5480
rect 25773 5475 25839 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 26532 5448 27332 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 25773 4858 25839 4861
rect 26532 4858 27332 4888
rect 25773 4856 27332 4858
rect 25773 4800 25778 4856
rect 25834 4800 27332 4856
rect 25773 4798 27332 4800
rect 25773 4795 25839 4798
rect 26532 4768 27332 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 20161 4178 20227 4181
rect 20529 4178 20595 4181
rect 20161 4176 20595 4178
rect 20161 4120 20166 4176
rect 20222 4120 20534 4176
rect 20590 4120 20595 4176
rect 20161 4118 20595 4120
rect 20161 4115 20227 4118
rect 20529 4115 20595 4118
rect 25405 4178 25471 4181
rect 26532 4178 27332 4208
rect 25405 4176 27332 4178
rect 25405 4120 25410 4176
rect 25466 4120 27332 4176
rect 25405 4118 27332 4120
rect 25405 4115 25471 4118
rect 26532 4088 27332 4118
rect 17493 4042 17559 4045
rect 23473 4042 23539 4045
rect 17493 4040 23539 4042
rect 17493 3984 17498 4040
rect 17554 3984 23478 4040
rect 23534 3984 23539 4040
rect 17493 3982 23539 3984
rect 17493 3979 17559 3982
rect 23473 3979 23539 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 19701 3636 19767 3637
rect 19701 3632 19748 3636
rect 19812 3634 19818 3636
rect 20529 3634 20595 3637
rect 23841 3634 23907 3637
rect 19701 3576 19706 3632
rect 19701 3572 19748 3576
rect 19812 3574 19858 3634
rect 20529 3632 23907 3634
rect 20529 3576 20534 3632
rect 20590 3576 23846 3632
rect 23902 3576 23907 3632
rect 20529 3574 23907 3576
rect 19812 3572 19818 3574
rect 19701 3571 19767 3572
rect 20529 3571 20595 3574
rect 23841 3571 23907 3574
rect 25773 3498 25839 3501
rect 26532 3498 27332 3528
rect 25773 3496 27332 3498
rect 25773 3440 25778 3496
rect 25834 3440 27332 3496
rect 25773 3438 27332 3440
rect 25773 3435 25839 3438
rect 26532 3408 27332 3438
rect 19425 3362 19491 3365
rect 20897 3362 20963 3365
rect 19425 3360 20963 3362
rect 19425 3304 19430 3360
rect 19486 3304 20902 3360
rect 20958 3304 20963 3360
rect 19425 3302 20963 3304
rect 19425 3299 19491 3302
rect 20897 3299 20963 3302
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 19701 3228 19767 3229
rect 19701 3226 19748 3228
rect 19656 3224 19748 3226
rect 19656 3168 19706 3224
rect 19656 3166 19748 3168
rect 19701 3164 19748 3166
rect 19812 3164 19818 3228
rect 20161 3226 20227 3229
rect 21449 3226 21515 3229
rect 20161 3224 21515 3226
rect 20161 3168 20166 3224
rect 20222 3168 21454 3224
rect 21510 3168 21515 3224
rect 20161 3166 21515 3168
rect 19701 3163 19767 3164
rect 20161 3163 20227 3166
rect 21449 3163 21515 3166
rect 16941 3090 17007 3093
rect 17125 3090 17191 3093
rect 22093 3090 22159 3093
rect 16941 3088 22159 3090
rect 16941 3032 16946 3088
rect 17002 3032 17130 3088
rect 17186 3032 22098 3088
rect 22154 3032 22159 3088
rect 16941 3030 22159 3032
rect 16941 3027 17007 3030
rect 17125 3027 17191 3030
rect 22093 3027 22159 3030
rect 20621 2954 20687 2957
rect 21081 2954 21147 2957
rect 20621 2952 21147 2954
rect 20621 2896 20626 2952
rect 20682 2896 21086 2952
rect 21142 2896 21147 2952
rect 20621 2894 21147 2896
rect 20621 2891 20687 2894
rect 21081 2891 21147 2894
rect 25773 2818 25839 2821
rect 26532 2818 27332 2848
rect 25773 2816 27332 2818
rect 25773 2760 25778 2816
rect 25834 2760 27332 2816
rect 25773 2758 27332 2760
rect 25773 2755 25839 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 26532 2728 27332 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 13492 23488 13556 23492
rect 13492 23432 13542 23488
rect 13542 23432 13556 23488
rect 13492 23428 13556 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 21220 23080 21284 23084
rect 21220 23024 21234 23080
rect 21234 23024 21284 23080
rect 21220 23020 21284 23024
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 21956 20768 22020 20772
rect 21956 20712 22006 20768
rect 22006 20712 22020 20768
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 21956 20708 22020 20712
rect 21220 20572 21284 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4660 19212 4724 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 13492 18456 13556 18460
rect 13492 18400 13542 18456
rect 13542 18400 13556 18456
rect 13492 18396 13556 18400
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 21956 15600 22020 15604
rect 21956 15544 21970 15600
rect 21970 15544 22020 15600
rect 21956 15540 22020 15544
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4660 11732 4724 11796
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 19748 3632 19812 3636
rect 19748 3576 19762 3632
rect 19762 3576 19812 3632
rect 19748 3572 19812 3576
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 19748 3224 19812 3228
rect 19748 3168 19762 3224
rect 19762 3168 19812 3224
rect 19748 3164 19812 3168
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 26688 4528 27248
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4868 27232 5188 27248
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4659 19276 4725 19277
rect 4659 19212 4660 19276
rect 4724 19212 4725 19276
rect 4659 19211 4725 19212
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4662 11797 4722 19211
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 13494 18461 13554 23427
rect 21219 23084 21285 23085
rect 21219 23020 21220 23084
rect 21284 23020 21285 23084
rect 21219 23019 21285 23020
rect 21222 20637 21282 23019
rect 21955 20772 22021 20773
rect 21955 20708 21956 20772
rect 22020 20708 22021 20772
rect 21955 20707 22021 20708
rect 21219 20636 21285 20637
rect 21219 20572 21220 20636
rect 21284 20572 21285 20636
rect 21219 20571 21285 20572
rect 13491 18460 13557 18461
rect 13491 18396 13492 18460
rect 13556 18396 13557 18460
rect 13491 18395 13557 18396
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 21958 15605 22018 20707
rect 21955 15604 22021 15605
rect 21955 15540 21956 15604
rect 22020 15540 22021 15604
rect 21955 15539 22021 15540
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4659 11796 4725 11797
rect 4659 11732 4660 11796
rect 4724 11732 4725 11796
rect 4659 11731 4725 11732
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 19747 3636 19813 3637
rect 19747 3572 19748 3636
rect 19812 3572 19813 3636
rect 19747 3571 19813 3572
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 19750 3229 19810 3571
rect 19747 3228 19813 3229
rect 19747 3164 19748 3228
rect 19812 3164 19813 3228
rect 19747 3163 19813 3164
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0527_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 11776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1730889744
transform -1 0 20148 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1730889744
transform 1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1730889744
transform -1 0 19044 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1730889744
transform -1 0 17756 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1730889744
transform 1 0 17848 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1730889744
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1730889744
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1730889744
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1730889744
transform 1 0 20056 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1730889744
transform 1 0 4508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0538_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0539_
timestamp 1730889744
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0540_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 11776 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0541_
timestamp 1730889744
transform 1 0 12420 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0542_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 13892 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0543_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 12788 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0544_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 13432 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0545_
timestamp 1730889744
transform 1 0 10396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0546_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10764 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1730889744
transform 1 0 6348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1730889744
transform -1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0549_
timestamp 1730889744
transform -1 0 8556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0550_
timestamp 1730889744
transform 1 0 7636 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0551_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5704 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0552_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 6808 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0553_
timestamp 1730889744
transform 1 0 6624 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0554_
timestamp 1730889744
transform -1 0 8188 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0555_
timestamp 1730889744
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0556_
timestamp 1730889744
transform 1 0 4232 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0557_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5244 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _0558_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 2944 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0559_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 5796 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0560_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0561_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0562_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5888 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0563_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 4048 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1730889744
transform 1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0565_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0566_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 5428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0567_
timestamp 1730889744
transform -1 0 5796 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0568_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 5244 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0569_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5244 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0570_
timestamp 1730889744
transform -1 0 5428 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0571_
timestamp 1730889744
transform -1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0572_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 6072 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0573_
timestamp 1730889744
transform -1 0 5428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0574_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5152 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0575_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 6164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0576_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 7452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0577_
timestamp 1730889744
transform 1 0 8188 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0578_
timestamp 1730889744
transform -1 0 8372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0579_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 7636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _0580_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 6348 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0581_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0582_
timestamp 1730889744
transform 1 0 6348 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _0583_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 7084 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0584_
timestamp 1730889744
transform 1 0 10028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0585_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 13248 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1730889744
transform 1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0587_
timestamp 1730889744
transform 1 0 14812 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0588_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 15364 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _0589_
timestamp 1730889744
transform 1 0 11776 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _0590_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 11776 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _0591_
timestamp 1730889744
transform -1 0 16560 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0592_
timestamp 1730889744
transform 1 0 16928 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0593_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 21620 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0594_
timestamp 1730889744
transform -1 0 21620 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0595_
timestamp 1730889744
transform -1 0 22172 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0596_
timestamp 1730889744
transform 1 0 20884 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1730889744
transform 1 0 21160 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0598_
timestamp 1730889744
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0599_
timestamp 1730889744
transform 1 0 23276 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0600_
timestamp 1730889744
transform -1 0 22632 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0601_
timestamp 1730889744
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0602_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 11960 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0603_
timestamp 1730889744
transform 1 0 11316 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0604_
timestamp 1730889744
transform 1 0 17480 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0605_
timestamp 1730889744
transform 1 0 20332 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0606_
timestamp 1730889744
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0607_
timestamp 1730889744
transform 1 0 18676 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0608_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 19688 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0609_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 19320 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0610_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0611_
timestamp 1730889744
transform 1 0 22540 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1730889744
transform 1 0 22632 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1730889744
transform -1 0 24748 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0614_
timestamp 1730889744
transform 1 0 7544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0615_
timestamp 1730889744
transform 1 0 7544 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0616_
timestamp 1730889744
transform 1 0 6716 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0617_
timestamp 1730889744
transform 1 0 7360 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0618_
timestamp 1730889744
transform 1 0 3956 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0619_
timestamp 1730889744
transform -1 0 4140 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0620_
timestamp 1730889744
transform 1 0 4416 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0621_
timestamp 1730889744
transform 1 0 5612 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0622_
timestamp 1730889744
transform -1 0 5612 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1730889744
transform -1 0 7268 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0624_
timestamp 1730889744
transform -1 0 6532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1730889744
transform 1 0 4232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0626_
timestamp 1730889744
transform 1 0 3588 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0627_
timestamp 1730889744
transform 1 0 5520 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0628_
timestamp 1730889744
transform 1 0 6532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0629_
timestamp 1730889744
transform 1 0 4232 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0630_
timestamp 1730889744
transform -1 0 5060 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0631_
timestamp 1730889744
transform 1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0632_
timestamp 1730889744
transform -1 0 5152 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0633_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 5336 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0634_
timestamp 1730889744
transform -1 0 5888 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0635_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0636_
timestamp 1730889744
transform -1 0 6900 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1730889744
transform -1 0 6716 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0638_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 7544 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _0639_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 6716 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0640_
timestamp 1730889744
transform 1 0 5428 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0641_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0642_
timestamp 1730889744
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0643_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 2852 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1730889744
transform 1 0 2024 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0645_
timestamp 1730889744
transform -1 0 3588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0646_
timestamp 1730889744
transform -1 0 3220 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0647_
timestamp 1730889744
transform -1 0 3036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1730889744
transform -1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0649_
timestamp 1730889744
transform -1 0 2760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0650_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 3220 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1730889744
transform 1 0 3312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0652_
timestamp 1730889744
transform 1 0 3496 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0653_
timestamp 1730889744
transform -1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0654_
timestamp 1730889744
transform -1 0 3864 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0655_
timestamp 1730889744
transform -1 0 3220 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0656_
timestamp 1730889744
transform 1 0 4140 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1730889744
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1730889744
transform -1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0659_
timestamp 1730889744
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1730889744
transform 1 0 5244 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1730889744
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1730889744
transform -1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0663_
timestamp 1730889744
transform 1 0 4876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0664_
timestamp 1730889744
transform 1 0 6348 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0665_
timestamp 1730889744
transform -1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0666_
timestamp 1730889744
transform 1 0 7176 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0667_
timestamp 1730889744
transform -1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1730889744
transform 1 0 8280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0669_
timestamp 1730889744
transform 1 0 7544 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1730889744
transform -1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1730889744
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0672_
timestamp 1730889744
transform -1 0 8740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0673_
timestamp 1730889744
transform 1 0 7728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1730889744
transform -1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0675_
timestamp 1730889744
transform 1 0 8188 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0676_
timestamp 1730889744
transform -1 0 10856 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1730889744
transform -1 0 8924 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0678_
timestamp 1730889744
transform 1 0 7912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0679_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 8832 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0680_
timestamp 1730889744
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0681_
timestamp 1730889744
transform 1 0 10672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0682_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0683_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 11592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1730889744
transform -1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 1730889744
transform 1 0 12420 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0686_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 12420 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1730889744
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0688_
timestamp 1730889744
transform 1 0 17756 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0689_
timestamp 1730889744
transform -1 0 17756 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0690_
timestamp 1730889744
transform -1 0 13984 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0691_
timestamp 1730889744
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1730889744
transform 1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0693_
timestamp 1730889744
transform -1 0 21252 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0694_
timestamp 1730889744
transform -1 0 21620 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1730889744
transform 1 0 19964 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1730889744
transform -1 0 14444 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0697_
timestamp 1730889744
transform 1 0 13248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0698_
timestamp 1730889744
transform -1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0699_
timestamp 1730889744
transform -1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0700_
timestamp 1730889744
transform 1 0 14076 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0701_
timestamp 1730889744
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0702_
timestamp 1730889744
transform -1 0 21712 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0703_
timestamp 1730889744
transform 1 0 20148 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1730889744
transform -1 0 17204 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0705_
timestamp 1730889744
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0706_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1730889744
transform 1 0 22172 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0708_
timestamp 1730889744
transform -1 0 21712 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0709_
timestamp 1730889744
transform 1 0 25300 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1730889744
transform -1 0 23828 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0711_
timestamp 1730889744
transform -1 0 24840 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0712_
timestamp 1730889744
transform -1 0 24288 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0713_
timestamp 1730889744
transform -1 0 25300 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0714_
timestamp 1730889744
transform -1 0 24104 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1730889744
transform -1 0 25300 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0716_
timestamp 1730889744
transform -1 0 23920 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0717_
timestamp 1730889744
transform 1 0 23828 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0718_
timestamp 1730889744
transform -1 0 25116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0719_
timestamp 1730889744
transform -1 0 23920 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0720_
timestamp 1730889744
transform -1 0 23920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1730889744
transform -1 0 22908 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0722_
timestamp 1730889744
transform 1 0 21712 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1730889744
transform -1 0 23000 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0724_
timestamp 1730889744
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _0725_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 19964 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1730889744
transform 1 0 21160 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0727_
timestamp 1730889744
transform 1 0 20240 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1730889744
transform 1 0 25024 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0729_
timestamp 1730889744
transform -1 0 24288 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1730889744
transform 1 0 24104 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0731_
timestamp 1730889744
transform -1 0 25116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0732_
timestamp 1730889744
transform -1 0 24104 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0733_
timestamp 1730889744
transform 1 0 22632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1730889744
transform -1 0 23828 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0735_
timestamp 1730889744
transform -1 0 24104 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0736_
timestamp 1730889744
transform 1 0 21252 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0737_
timestamp 1730889744
transform -1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1730889744
transform -1 0 24288 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0739_
timestamp 1730889744
transform -1 0 23644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0740_
timestamp 1730889744
transform 1 0 21160 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0741_
timestamp 1730889744
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0742_
timestamp 1730889744
transform 1 0 21252 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0743_
timestamp 1730889744
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0744_
timestamp 1730889744
transform -1 0 18768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1730889744
transform -1 0 18492 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0746_
timestamp 1730889744
transform 1 0 17572 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1730889744
transform -1 0 16100 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1730889744
transform 1 0 14352 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1730889744
transform -1 0 17940 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0750_
timestamp 1730889744
transform -1 0 17848 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1730889744
transform 1 0 19412 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0752_
timestamp 1730889744
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1730889744
transform -1 0 15640 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1730889744
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1730889744
transform 1 0 18400 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1730889744
transform 1 0 19596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1730889744
transform -1 0 17480 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1730889744
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1730889744
transform 1 0 16652 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1730889744
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1730889744
transform -1 0 19688 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1730889744
transform 1 0 18032 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0763_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1730889744
transform 1 0 18676 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0765_
timestamp 1730889744
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0766_
timestamp 1730889744
transform -1 0 18400 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0767_
timestamp 1730889744
transform -1 0 19136 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1730889744
transform 1 0 23092 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0769_
timestamp 1730889744
transform -1 0 24288 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1730889744
transform 1 0 24380 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0771_
timestamp 1730889744
transform -1 0 23828 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1730889744
transform 1 0 20332 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0773_
timestamp 1730889744
transform -1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1730889744
transform 1 0 24380 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0775_
timestamp 1730889744
transform -1 0 24380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1730889744
transform -1 0 20056 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0777_
timestamp 1730889744
transform 1 0 18860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1730889744
transform -1 0 22264 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0779_
timestamp 1730889744
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1730889744
transform -1 0 23092 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0781_
timestamp 1730889744
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1730889744
transform -1 0 16468 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1730889744
transform -1 0 25024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0784_
timestamp 1730889744
transform 1 0 14996 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1730889744
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1730889744
transform 1 0 19964 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1730889744
transform -1 0 24012 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0788_
timestamp 1730889744
transform 1 0 19872 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1730889744
transform 1 0 17848 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0790_
timestamp 1730889744
transform 1 0 20332 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0791_
timestamp 1730889744
transform -1 0 25024 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0792_
timestamp 1730889744
transform 1 0 20700 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1730889744
transform 1 0 18492 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1730889744
transform -1 0 25760 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0795_
timestamp 1730889744
transform -1 0 16468 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0796_
timestamp 1730889744
transform 1 0 14904 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1730889744
transform -1 0 15640 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1730889744
transform -1 0 25760 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1730889744
transform -1 0 20884 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0800_
timestamp 1730889744
transform 1 0 19504 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1730889744
transform 1 0 18584 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0802_
timestamp 1730889744
transform -1 0 17296 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0803_
timestamp 1730889744
transform -1 0 25024 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0804_
timestamp 1730889744
transform 1 0 14904 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1730889744
transform -1 0 13984 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1730889744
transform -1 0 22632 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1730889744
transform 1 0 20884 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0808_
timestamp 1730889744
transform 1 0 20516 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1730889744
transform 1 0 19412 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1730889744
transform -1 0 20608 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1730889744
transform -1 0 22448 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0812_
timestamp 1730889744
transform 1 0 16652 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1730889744
transform 1 0 16652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1730889744
transform 1 0 17940 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1730889744
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1730889744
transform 1 0 17296 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0817_
timestamp 1730889744
transform 1 0 14628 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1730889744
transform 1 0 15364 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0819_
timestamp 1730889744
transform 1 0 14536 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1730889744
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0821_
timestamp 1730889744
transform -1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1730889744
transform 1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1730889744
transform -1 0 13984 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1730889744
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0825_
timestamp 1730889744
transform 1 0 13248 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0826_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10488 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1730889744
transform -1 0 11868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1730889744
transform 1 0 11960 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1730889744
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1730889744
transform -1 0 14444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1730889744
transform 1 0 11500 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0832_
timestamp 1730889744
transform 1 0 12052 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1730889744
transform 1 0 11868 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1730889744
transform 1 0 12420 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1730889744
transform 1 0 14996 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1730889744
transform 1 0 12052 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0837_
timestamp 1730889744
transform -1 0 14444 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0838_
timestamp 1730889744
transform 1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0839_
timestamp 1730889744
transform -1 0 13984 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0840_
timestamp 1730889744
transform 1 0 12512 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1730889744
transform -1 0 13984 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1730889744
transform 1 0 13984 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1730889744
transform -1 0 13616 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0844_
timestamp 1730889744
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0845_
timestamp 1730889744
transform 1 0 12236 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1730889744
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0847_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10856 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1730889744
transform 1 0 11868 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1730889744
transform 1 0 16652 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1730889744
transform 1 0 14812 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1730889744
transform 1 0 17388 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1730889744
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1730889744
transform 1 0 14444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1730889744
transform 1 0 12420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1730889744
transform 1 0 18216 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1730889744
transform 1 0 12972 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1730889744
transform -1 0 16284 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1730889744
transform 1 0 15548 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1730889744
transform 1 0 17848 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1730889744
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1730889744
transform 1 0 17848 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1730889744
transform -1 0 15824 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1730889744
transform 1 0 15180 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1730889744
transform -1 0 14996 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1730889744
transform 1 0 6256 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1730889744
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0867_
timestamp 1730889744
transform -1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1730889744
transform -1 0 4784 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0869_
timestamp 1730889744
transform -1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1730889744
transform -1 0 3680 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1730889744
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0872_
timestamp 1730889744
transform 1 0 4784 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1730889744
transform 1 0 8740 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1730889744
transform 1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1730889744
transform 1 0 6900 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 1730889744
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_1  _0877_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 7452 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0878_
timestamp 1730889744
transform -1 0 8740 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0879_
timestamp 1730889744
transform -1 0 8096 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0880_
timestamp 1730889744
transform -1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1730889744
transform 1 0 2852 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1730889744
transform -1 0 4692 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0883_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0884_
timestamp 1730889744
transform -1 0 2760 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0885_
timestamp 1730889744
transform 1 0 3772 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0886_
timestamp 1730889744
transform 1 0 2760 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0887_
timestamp 1730889744
transform -1 0 2852 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1730889744
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0889_
timestamp 1730889744
transform -1 0 2208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1730889744
transform -1 0 3588 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1730889744
transform -1 0 4324 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1730889744
transform 1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0893_
timestamp 1730889744
transform 1 0 2208 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0894_
timestamp 1730889744
transform -1 0 5704 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1730889744
transform 1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0896_
timestamp 1730889744
transform -1 0 6256 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1730889744
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1730889744
transform -1 0 5244 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1730889744
transform 1 0 5152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0900_
timestamp 1730889744
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1730889744
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0902_
timestamp 1730889744
transform -1 0 6164 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1730889744
transform 1 0 7268 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1730889744
transform 1 0 7452 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0905_
timestamp 1730889744
transform 1 0 8188 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1730889744
transform -1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1730889744
transform 1 0 9016 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1730889744
transform -1 0 9936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0909_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 7728 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1730889744
transform -1 0 12420 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1730889744
transform -1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1730889744
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1730889744
transform -1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0914_
timestamp 1730889744
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1730889744
transform -1 0 13984 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0916_
timestamp 1730889744
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0917_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1730889744
transform 1 0 11316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0919_
timestamp 1730889744
transform -1 0 13984 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1730889744
transform -1 0 12880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0921_
timestamp 1730889744
transform 1 0 12972 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0922_
timestamp 1730889744
transform -1 0 11960 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1730889744
transform -1 0 11408 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0924_
timestamp 1730889744
transform 1 0 10212 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1730889744
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0926_
timestamp 1730889744
transform -1 0 2392 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1730889744
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1730889744
transform -1 0 3588 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1730889744
transform 1 0 2392 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1730889744
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1730889744
transform -1 0 3680 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1730889744
transform -1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0933_
timestamp 1730889744
transform -1 0 2852 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0934_
timestamp 1730889744
transform -1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1730889744
transform 1 0 3036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1730889744
transform 1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1730889744
transform -1 0 2576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1730889744
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1730889744
transform -1 0 3220 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0940_
timestamp 1730889744
transform -1 0 2760 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0941_
timestamp 1730889744
transform -1 0 3588 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0942_
timestamp 1730889744
transform -1 0 4600 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1730889744
transform -1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1730889744
transform -1 0 3680 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0945_
timestamp 1730889744
transform 1 0 3588 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1730889744
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1730889744
transform 1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1730889744
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0949_
timestamp 1730889744
transform 1 0 4692 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1730889744
transform -1 0 5888 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1730889744
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1730889744
transform -1 0 7176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1730889744
transform 1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0954_
timestamp 1730889744
transform 1 0 7176 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0955_
timestamp 1730889744
transform 1 0 7636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1730889744
transform 1 0 8280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1730889744
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0958_
timestamp 1730889744
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0959_
timestamp 1730889744
transform -1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1730889744
transform 1 0 8740 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0961_
timestamp 1730889744
transform -1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1730889744
transform 1 0 9384 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1730889744
transform 1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0964_
timestamp 1730889744
transform 1 0 8372 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1730889744
transform -1 0 9384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0966_
timestamp 1730889744
transform 1 0 21804 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0967_
timestamp 1730889744
transform -1 0 23092 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0968_
timestamp 1730889744
transform 1 0 23552 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1730889744
transform 1 0 24380 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1730889744
transform 1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1730889744
transform 1 0 12880 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1730889744
transform 1 0 19872 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1730889744
transform 1 0 19688 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0974_
timestamp 1730889744
transform 1 0 18768 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0975_
timestamp 1730889744
transform -1 0 18768 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0976_
timestamp 1730889744
transform -1 0 21436 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0977_
timestamp 1730889744
transform 1 0 20976 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1730889744
transform 1 0 20424 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0979_
timestamp 1730889744
transform 1 0 20608 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0980_
timestamp 1730889744
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0981_
timestamp 1730889744
transform 1 0 19964 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1730889744
transform -1 0 20240 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1730889744
transform 1 0 19412 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1730889744
transform -1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0985_
timestamp 1730889744
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1730889744
transform 1 0 20240 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0987_
timestamp 1730889744
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1730889744
transform -1 0 20976 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1730889744
transform -1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0990_
timestamp 1730889744
transform 1 0 18308 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1730889744
transform -1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1730889744
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0993_
timestamp 1730889744
transform 1 0 20884 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0994_
timestamp 1730889744
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0995_
timestamp 1730889744
transform 1 0 21620 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0996_
timestamp 1730889744
transform -1 0 22172 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0997_
timestamp 1730889744
transform -1 0 21528 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1730889744
transform 1 0 18676 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0999_
timestamp 1730889744
transform 1 0 21436 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1000_
timestamp 1730889744
transform -1 0 18860 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1730889744
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1002_
timestamp 1730889744
transform -1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1730889744
transform 1 0 22080 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1730889744
transform 1 0 22816 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1730889744
transform 1 0 24380 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1006_
timestamp 1730889744
transform 1 0 20792 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1007_
timestamp 1730889744
transform -1 0 22172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1008_
timestamp 1730889744
transform 1 0 23276 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1730889744
transform -1 0 24288 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 1730889744
transform 1 0 21804 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1730889744
transform -1 0 22540 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1012_
timestamp 1730889744
transform -1 0 23552 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1013_
timestamp 1730889744
transform 1 0 23092 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1730889744
transform 1 0 24380 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1015_
timestamp 1730889744
transform 1 0 21620 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1016_
timestamp 1730889744
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 1730889744
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1730889744
transform 1 0 22264 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1730889744
transform -1 0 24288 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1020_
timestamp 1730889744
transform -1 0 20332 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1021_
timestamp 1730889744
transform 1 0 20332 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1022_
timestamp 1730889744
transform -1 0 20332 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1023_
timestamp 1730889744
transform 1 0 20332 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1024_
timestamp 1730889744
transform 1 0 21620 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1730889744
transform -1 0 22356 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1730889744
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1027_
timestamp 1730889744
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1730889744
transform -1 0 21436 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1029_
timestamp 1730889744
transform -1 0 21160 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1030_
timestamp 1730889744
transform 1 0 19228 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 1730889744
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1730889744
transform -1 0 12328 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1033_
timestamp 1730889744
transform 1 0 12420 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1034_
timestamp 1730889744
transform -1 0 13340 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1730889744
transform -1 0 12512 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1730889744
transform -1 0 12420 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1730889744
transform -1 0 20240 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1730889744
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1730889744
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1040_
timestamp 1730889744
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 1730889744
transform 1 0 14076 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1042_
timestamp 1730889744
transform 1 0 14168 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 1730889744
transform 1 0 15640 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1044_
timestamp 1730889744
transform 1 0 16744 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1730889744
transform 1 0 18768 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1730889744
transform -1 0 16560 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1047_
timestamp 1730889744
transform 1 0 18216 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1730889744
transform -1 0 13984 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1049_
timestamp 1730889744
transform 1 0 13248 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1730889744
transform -1 0 14720 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1730889744
transform -1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1730889744
transform -1 0 18768 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1053_
timestamp 1730889744
transform 1 0 20792 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1730889744
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1055_
timestamp 1730889744
transform 1 0 22908 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 1730889744
transform 1 0 24380 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1057_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 15272 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1058_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 24380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1730889744
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1730889744
transform -1 0 3312 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1730889744
transform 1 0 1840 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1730889744
transform 1 0 2024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1730889744
transform 1 0 2208 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1730889744
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1730889744
transform 1 0 4968 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1730889744
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1730889744
transform 1 0 7636 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1730889744
transform -1 0 8832 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1730889744
transform -1 0 10120 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1730889744
transform -1 0 10396 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1730889744
transform -1 0 10396 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1730889744
transform 1 0 10488 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1730889744
transform -1 0 13708 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1730889744
transform 1 0 12604 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1730889744
transform 1 0 20884 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1730889744
transform 1 0 19596 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1730889744
transform 1 0 12512 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1730889744
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1730889744
transform 1 0 13248 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1730889744
transform 1 0 20240 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1730889744
transform 1 0 15088 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1730889744
transform 1 0 23828 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1730889744
transform 1 0 23828 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1730889744
transform 1 0 24104 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1730889744
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1730889744
transform 1 0 24012 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1730889744
transform 1 0 24380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1730889744
transform 1 0 21804 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1730889744
transform 1 0 21068 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1730889744
transform 1 0 24380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1730889744
transform -1 0 24932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1730889744
transform 1 0 22632 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1730889744
transform 1 0 24104 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1730889744
transform 1 0 22172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1730889744
transform 1 0 23644 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1730889744
transform -1 0 22172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1730889744
transform 1 0 21804 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1730889744
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1730889744
transform 1 0 17296 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1730889744
transform 1 0 18124 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1730889744
transform 1 0 13708 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1730889744
transform -1 0 19412 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1730889744
transform 1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1730889744
transform 1 0 15824 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1730889744
transform 1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1730889744
transform 1 0 19228 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1730889744
transform 1 0 24380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1730889744
transform 1 0 23828 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1730889744
transform 1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1730889744
transform 1 0 24380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1730889744
transform 1 0 19044 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1730889744
transform 1 0 20884 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1730889744
transform 1 0 20700 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1730889744
transform 1 0 13524 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1730889744
transform -1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1730889744
transform 1 0 17112 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1730889744
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1730889744
transform 1 0 15088 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1730889744
transform 1 0 17388 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1730889744
transform 1 0 13708 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1730889744
transform 1 0 17112 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1730889744
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1730889744
transform 1 0 17572 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1730889744
transform 1 0 17572 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1730889744
transform 1 0 17020 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1126_
timestamp 1730889744
transform 1 0 14996 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1127_
timestamp 1730889744
transform 1 0 15180 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1730889744
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1730889744
transform -1 0 10856 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1730889744
transform 1 0 11776 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1730889744
transform 1 0 11500 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1730889744
transform 1 0 12512 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1730889744
transform -1 0 15640 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1730889744
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1730889744
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1730889744
transform -1 0 12420 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1730889744
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1730889744
transform -1 0 15548 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1730889744
transform -1 0 15916 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1730889744
transform -1 0 14996 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1730889744
transform 1 0 2116 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1730889744
transform -1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1730889744
transform 1 0 1932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1730889744
transform 1 0 2024 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1730889744
transform -1 0 3128 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1730889744
transform 1 0 2852 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1730889744
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1730889744
transform -1 0 8188 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1730889744
transform 1 0 5244 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1730889744
transform -1 0 9384 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1730889744
transform -1 0 10396 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1730889744
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1730889744
transform 1 0 9936 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1730889744
transform 1 0 8188 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1730889744
transform 1 0 9292 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1730889744
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1730889744
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1730889744
transform -1 0 12972 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1730889744
transform 1 0 12052 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1730889744
transform 1 0 9844 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1730889744
transform 1 0 9936 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1730889744
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1730889744
transform 1 0 11040 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1730889744
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1730889744
transform 1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1730889744
transform 1 0 2300 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1730889744
transform 1 0 1748 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1730889744
transform 1 0 1656 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1730889744
transform 1 0 2024 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1730889744
transform -1 0 4324 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1730889744
transform 1 0 5336 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1730889744
transform -1 0 9016 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1730889744
transform -1 0 9752 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1730889744
transform -1 0 10672 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1730889744
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1730889744
transform -1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1730889744
transform 1 0 23736 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1178_
timestamp 1730889744
transform 1 0 11316 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1730889744
transform -1 0 18124 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1730889744
transform -1 0 18952 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1730889744
transform 1 0 16928 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1730889744
transform -1 0 18308 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1730889744
transform -1 0 20056 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1730889744
transform -1 0 21712 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1730889744
transform 1 0 16928 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1730889744
transform 1 0 23368 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1730889744
transform 1 0 23736 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1730889744
transform 1 0 23828 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1730889744
transform 1 0 24380 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1730889744
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1730889744
transform 1 0 22816 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1730889744
transform -1 0 23092 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1730889744
transform -1 0 21620 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1730889744
transform 1 0 19044 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1730889744
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1730889744
transform 1 0 11684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1730889744
transform 1 0 11500 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1730889744
transform 1 0 15640 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1730889744
transform -1 0 15732 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1200_
timestamp 1730889744
transform 1 0 13800 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1201_
timestamp 1730889744
transform 1 0 14720 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1730889744
transform 1 0 16468 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1730889744
transform -1 0 18216 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1204_
timestamp 1730889744
transform 1 0 14076 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1205_
timestamp 1730889744
transform 1 0 14076 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1730889744
transform -1 0 18124 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1730889744
transform 1 0 23736 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1208_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1730889744
transform -1 0 23736 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1730889744
transform -1 0 23828 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1730889744
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1730889744
transform 1 0 25300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1730889744
transform -1 0 25484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1730889744
transform -1 0 25024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1730889744
transform -1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 13248 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 4048 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1730889744
transform -1 0 4784 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1730889744
transform 1 0 9660 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1730889744
transform 1 0 10212 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1730889744
transform -1 0 6256 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1730889744
transform -1 0 9568 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1730889744
transform 1 0 11040 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1730889744
transform 1 0 10488 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1730889744
transform -1 0 16744 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1730889744
transform 1 0 16652 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1730889744
transform 1 0 21804 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1730889744
transform 1 0 22172 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1730889744
transform 1 0 16836 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1730889744
transform 1 0 17204 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1730889744
transform 1 0 22264 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1730889744
transform 1 0 22264 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 4048 0 -1 9792
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 3680 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp 1730889744
transform 1 0 10764 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload3
timestamp 1730889744
transform 1 0 10212 0 1 9792
box -38 -48 2246 592
use sky130_fd_sc_hd__bufinv_16  clkload4
timestamp 1730889744
transform 1 0 6348 0 -1 20672
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  clkload5 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 9568 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  clkload6 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10488 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload7
timestamp 1730889744
transform 1 0 11500 0 1 19584
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload8
timestamp 1730889744
transform -1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload9
timestamp 1730889744
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload10
timestamp 1730889744
transform 1 0 22448 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload11
timestamp 1730889744
transform 1 0 16836 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload12
timestamp 1730889744
transform 1 0 22264 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__bufinv_16  clkload13
timestamp 1730889744
transform 1 0 22080 0 1 17408
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_2  fanout58 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 6992 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1730889744
transform -1 0 9200 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1730889744
transform -1 0 10028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1730889744
transform -1 0 9660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout62
timestamp 1730889744
transform -1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1730889744
transform -1 0 13800 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout64 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform -1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 1730889744
transform -1 0 14536 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout67
timestamp 1730889744
transform -1 0 21436 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1730889744
transform -1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout69
timestamp 1730889744
transform 1 0 11040 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1730889744
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 1730889744
transform 1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 1730889744
transform -1 0 6716 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1730889744
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 1730889744
transform 1 0 21712 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1730889744
transform -1 0 19136 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1730889744
transform 1 0 21896 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout77
timestamp 1730889744
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 1730889744
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout79
timestamp 1730889744
transform -1 0 6808 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 1730889744
transform 1 0 4232 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout81
timestamp 1730889744
transform -1 0 4324 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1730889744
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1730889744
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1730889744
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1730889744
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1730889744
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1730889744
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1730889744
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1730889744
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp 1730889744
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1730889744
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_147
timestamp 1730889744
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp 1730889744
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp 1730889744
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1730889744
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp 1730889744
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1730889744
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1730889744
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1730889744
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_210
timestamp 1730889744
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1730889744
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1730889744
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1730889744
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_238
timestamp 1730889744
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_245
timestamp 1730889744
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1730889744
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_267
timestamp 1730889744
transform 1 0 25668 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1730889744
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1730889744
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1730889744
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1730889744
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1730889744
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1730889744
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1730889744
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1730889744
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1730889744
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1730889744
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1730889744
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1730889744
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1730889744
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1730889744
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1730889744
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1730889744
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1730889744
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1730889744
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1730889744
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1730889744
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp 1730889744
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_263
timestamp 1730889744
transform 1 0 25300 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1730889744
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1730889744
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1730889744
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1730889744
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1730889744
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1730889744
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1730889744
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1730889744
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1730889744
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1730889744
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1730889744
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1730889744
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1730889744
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1730889744
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1730889744
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_157
timestamp 1730889744
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_212
timestamp 1730889744
transform 1 0 20608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1730889744
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_261
timestamp 1730889744
transform 1 0 25116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_265
timestamp 1730889744
transform 1 0 25484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1730889744
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1730889744
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1730889744
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1730889744
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1730889744
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1730889744
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1730889744
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1730889744
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1730889744
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1730889744
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1730889744
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1730889744
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1730889744
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_141
timestamp 1730889744
transform 1 0 14076 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1730889744
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_182
timestamp 1730889744
transform 1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_216
timestamp 1730889744
transform 1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_233
timestamp 1730889744
transform 1 0 22540 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp 1730889744
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_259
timestamp 1730889744
transform 1 0 24932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1730889744
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1730889744
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1730889744
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1730889744
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1730889744
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1730889744
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1730889744
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1730889744
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1730889744
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1730889744
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_121
timestamp 1730889744
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_149
timestamp 1730889744
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1730889744
transform 1 0 15272 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_167
timestamp 1730889744
transform 1 0 16468 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1730889744
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1730889744
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_202
timestamp 1730889744
transform 1 0 19688 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1730889744
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_218
timestamp 1730889744
transform 1 0 21160 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_228
timestamp 1730889744
transform 1 0 22080 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1730889744
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_269
timestamp 1730889744
transform 1 0 25852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1730889744
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1730889744
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_47
timestamp 1730889744
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1730889744
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1730889744
transform 1 0 6808 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_68
timestamp 1730889744
transform 1 0 7360 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_90
timestamp 1730889744
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_102
timestamp 1730889744
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1730889744
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1730889744
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_125
timestamp 1730889744
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1730889744
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_145
timestamp 1730889744
transform 1 0 14444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1730889744
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1730889744
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1730889744
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_181
timestamp 1730889744
transform 1 0 17756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_201
timestamp 1730889744
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1730889744
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1730889744
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1730889744
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1730889744
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1730889744
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1730889744
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_37
timestamp 1730889744
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1730889744
transform 1 0 10396 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_118
timestamp 1730889744
transform 1 0 11960 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_130
timestamp 1730889744
transform 1 0 13064 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_134
timestamp 1730889744
transform 1 0 13432 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_149
timestamp 1730889744
transform 1 0 14812 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_178
timestamp 1730889744
transform 1 0 17480 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1730889744
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1730889744
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1730889744
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_205
timestamp 1730889744
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_229
timestamp 1730889744
transform 1 0 22172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_241
timestamp 1730889744
transform 1 0 23276 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1730889744
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1730889744
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_31
timestamp 1730889744
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1730889744
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1730889744
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_60
timestamp 1730889744
transform 1 0 6624 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1730889744
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_96
timestamp 1730889744
transform 1 0 9936 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1730889744
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_124
timestamp 1730889744
transform 1 0 12512 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_148
timestamp 1730889744
transform 1 0 14720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_156
timestamp 1730889744
transform 1 0 15456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1730889744
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_176
timestamp 1730889744
transform 1 0 17296 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_188
timestamp 1730889744
transform 1 0 18400 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_194
timestamp 1730889744
transform 1 0 18952 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_211
timestamp 1730889744
transform 1 0 20516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_217
timestamp 1730889744
transform 1 0 21068 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1730889744
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1730889744
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1730889744
transform 1 0 25760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1730889744
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1730889744
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_36
timestamp 1730889744
transform 1 0 4416 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_48
timestamp 1730889744
transform 1 0 5520 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1730889744
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_96
timestamp 1730889744
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_124
timestamp 1730889744
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1730889744
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1730889744
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1730889744
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_175
timestamp 1730889744
transform 1 0 17204 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp 1730889744
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_239
timestamp 1730889744
transform 1 0 23092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1730889744
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_260
timestamp 1730889744
transform 1 0 25024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1730889744
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1730889744
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1730889744
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40
timestamp 1730889744
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1730889744
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1730889744
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp 1730889744
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_88
timestamp 1730889744
transform 1 0 9200 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_100
timestamp 1730889744
transform 1 0 10304 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_127
timestamp 1730889744
transform 1 0 12788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_139
timestamp 1730889744
transform 1 0 13892 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1730889744
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_176
timestamp 1730889744
transform 1 0 17296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1730889744
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_192
timestamp 1730889744
transform 1 0 18768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_206
timestamp 1730889744
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1730889744
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1730889744
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1730889744
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1730889744
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1730889744
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1730889744
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_56
timestamp 1730889744
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1730889744
transform 1 0 7268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_101
timestamp 1730889744
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_110
timestamp 1730889744
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1730889744
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1730889744
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_173
timestamp 1730889744
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1730889744
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1730889744
transform 1 0 19688 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_210
timestamp 1730889744
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1730889744
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_269
timestamp 1730889744
transform 1 0 25852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1730889744
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_68
timestamp 1730889744
transform 1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_72
timestamp 1730889744
transform 1 0 7728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_155
timestamp 1730889744
transform 1 0 15364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1730889744
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_183
timestamp 1730889744
transform 1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_209
timestamp 1730889744
transform 1 0 20332 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1730889744
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_238
timestamp 1730889744
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_268
timestamp 1730889744
transform 1 0 25760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1730889744
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1730889744
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_67
timestamp 1730889744
transform 1 0 7268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1730889744
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1730889744
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1730889744
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1730889744
transform 1 0 14352 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1730889744
transform 1 0 15088 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_170
timestamp 1730889744
transform 1 0 16744 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_182
timestamp 1730889744
transform 1 0 17848 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_190
timestamp 1730889744
transform 1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1730889744
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_203
timestamp 1730889744
transform 1 0 19780 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1730889744
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1730889744
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_263
timestamp 1730889744
transform 1 0 25300 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1730889744
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1730889744
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1730889744
transform 1 0 3036 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1730889744
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1730889744
transform 1 0 3956 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1730889744
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1730889744
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_81
timestamp 1730889744
transform 1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_87
timestamp 1730889744
transform 1 0 9108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1730889744
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_150
timestamp 1730889744
transform 1 0 14904 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_178
timestamp 1730889744
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_203
timestamp 1730889744
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1730889744
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1730889744
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp 1730889744
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_230
timestamp 1730889744
transform 1 0 22264 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_238
timestamp 1730889744
transform 1 0 23000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_263
timestamp 1730889744
transform 1 0 25300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_269
timestamp 1730889744
transform 1 0 25852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1730889744
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1730889744
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 1730889744
transform 1 0 3036 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1730889744
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_52
timestamp 1730889744
transform 1 0 5888 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_64
timestamp 1730889744
transform 1 0 6992 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp 1730889744
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1730889744
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_96
timestamp 1730889744
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_123
timestamp 1730889744
transform 1 0 12420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1730889744
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_146
timestamp 1730889744
transform 1 0 14536 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1730889744
transform 1 0 15272 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_164
timestamp 1730889744
transform 1 0 16192 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_176
timestamp 1730889744
transform 1 0 17296 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1730889744
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_214
timestamp 1730889744
transform 1 0 20792 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_231
timestamp 1730889744
transform 1 0 22356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_243
timestamp 1730889744
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1730889744
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_260
timestamp 1730889744
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1730889744
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1730889744
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1730889744
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1730889744
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1730889744
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_67
timestamp 1730889744
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_86
timestamp 1730889744
transform 1 0 9016 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp 1730889744
transform 1 0 10120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1730889744
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1730889744
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_122
timestamp 1730889744
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_126
timestamp 1730889744
transform 1 0 12696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1730889744
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_142
timestamp 1730889744
transform 1 0 14168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1730889744
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1730889744
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1730889744
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1730889744
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_192
timestamp 1730889744
transform 1 0 18768 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_204
timestamp 1730889744
transform 1 0 19872 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_230
timestamp 1730889744
transform 1 0 22264 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1730889744
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1730889744
transform 1 0 1932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1730889744
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 1730889744
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1730889744
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1730889744
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1730889744
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_117
timestamp 1730889744
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1730889744
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1730889744
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1730889744
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1730889744
transform 1 0 16836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_175
timestamp 1730889744
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1730889744
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1730889744
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_237
timestamp 1730889744
transform 1 0 22908 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_243
timestamp 1730889744
transform 1 0 23460 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1730889744
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1730889744
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1730889744
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1730889744
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1730889744
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_94
timestamp 1730889744
transform 1 0 9752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1730889744
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1730889744
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1730889744
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_198
timestamp 1730889744
transform 1 0 19320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1730889744
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_241
timestamp 1730889744
transform 1 0 23276 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_263
timestamp 1730889744
transform 1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1730889744
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_32
timestamp 1730889744
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_48
timestamp 1730889744
transform 1 0 5520 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_60
timestamp 1730889744
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_72
timestamp 1730889744
transform 1 0 7728 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_92
timestamp 1730889744
transform 1 0 9568 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_104
timestamp 1730889744
transform 1 0 10672 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_110
timestamp 1730889744
transform 1 0 11224 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1730889744
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_167
timestamp 1730889744
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_175
timestamp 1730889744
transform 1 0 17204 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1730889744
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1730889744
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1730889744
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1730889744
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_234
timestamp 1730889744
transform 1 0 22632 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_246
timestamp 1730889744
transform 1 0 23736 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_268
timestamp 1730889744
transform 1 0 25760 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1730889744
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1730889744
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_22
timestamp 1730889744
transform 1 0 3128 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_34
timestamp 1730889744
transform 1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_42
timestamp 1730889744
transform 1 0 4968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1730889744
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1730889744
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1730889744
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1730889744
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1730889744
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1730889744
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1730889744
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1730889744
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1730889744
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1730889744
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1730889744
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1730889744
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_181
timestamp 1730889744
transform 1 0 17756 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_191
timestamp 1730889744
transform 1 0 18676 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_199
timestamp 1730889744
transform 1 0 19412 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1730889744
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1730889744
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1730889744
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1730889744
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1730889744
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1730889744
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_16
timestamp 1730889744
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1730889744
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1730889744
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_57
timestamp 1730889744
transform 1 0 6348 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_89
timestamp 1730889744
transform 1 0 9292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_101
timestamp 1730889744
transform 1 0 10396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_113
timestamp 1730889744
transform 1 0 11500 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_124
timestamp 1730889744
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1730889744
transform 1 0 13064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1730889744
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1730889744
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1730889744
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1730889744
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_236
timestamp 1730889744
transform 1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_269
timestamp 1730889744
transform 1 0 25852 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1730889744
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1730889744
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1730889744
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1730889744
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1730889744
transform 1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_98
timestamp 1730889744
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1730889744
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1730889744
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1730889744
transform 1 0 13156 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1730889744
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1730889744
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_241
timestamp 1730889744
transform 1 0 23276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1730889744
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1730889744
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_58
timestamp 1730889744
transform 1 0 6440 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1730889744
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_71
timestamp 1730889744
transform 1 0 7636 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_101
timestamp 1730889744
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1730889744
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1730889744
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1730889744
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1730889744
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_226
timestamp 1730889744
transform 1 0 21896 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_238
timestamp 1730889744
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1730889744
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 1730889744
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1730889744
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1730889744
transform 1 0 4784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1730889744
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_62
timestamp 1730889744
transform 1 0 6808 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_74
timestamp 1730889744
transform 1 0 7912 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1730889744
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1730889744
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_186
timestamp 1730889744
transform 1 0 18216 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_198
timestamp 1730889744
transform 1 0 19320 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_210
timestamp 1730889744
transform 1 0 20424 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1730889744
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1730889744
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_230
timestamp 1730889744
transform 1 0 22264 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_238
timestamp 1730889744
transform 1 0 23000 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_250
timestamp 1730889744
transform 1 0 24104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_258
timestamp 1730889744
transform 1 0 24840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_262
timestamp 1730889744
transform 1 0 25208 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1730889744
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1730889744
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_36
timestamp 1730889744
transform 1 0 4416 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_44
timestamp 1730889744
transform 1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_51
timestamp 1730889744
transform 1 0 5796 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1730889744
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1730889744
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1730889744
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1730889744
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_100
timestamp 1730889744
transform 1 0 10304 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1730889744
transform 1 0 10856 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1730889744
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1730889744
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_162
timestamp 1730889744
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_174
timestamp 1730889744
transform 1 0 17112 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1730889744
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1730889744
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1730889744
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_214
timestamp 1730889744
transform 1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_235
timestamp 1730889744
transform 1 0 22724 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_261
timestamp 1730889744
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_7
timestamp 1730889744
transform 1 0 1748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1730889744
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_39
timestamp 1730889744
transform 1 0 4692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1730889744
transform 1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1730889744
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_62
timestamp 1730889744
transform 1 0 6808 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_74
timestamp 1730889744
transform 1 0 7912 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_86
timestamp 1730889744
transform 1 0 9016 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_98
timestamp 1730889744
transform 1 0 10120 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1730889744
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_146
timestamp 1730889744
transform 1 0 14536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1730889744
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1730889744
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1730889744
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1730889744
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1730889744
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_228
timestamp 1730889744
transform 1 0 22080 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1730889744
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1730889744
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1730889744
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1730889744
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1730889744
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1730889744
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_67
timestamp 1730889744
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1730889744
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1730889744
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1730889744
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1730889744
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1730889744
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1730889744
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_125
timestamp 1730889744
transform 1 0 12604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1730889744
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1730889744
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_153
timestamp 1730889744
transform 1 0 15180 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_165
timestamp 1730889744
transform 1 0 16284 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_171
timestamp 1730889744
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1730889744
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1730889744
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1730889744
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_241
timestamp 1730889744
transform 1 0 23276 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 1730889744
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1730889744
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1730889744
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1730889744
transform 1 0 2852 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_27
timestamp 1730889744
transform 1 0 3588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_33
timestamp 1730889744
transform 1 0 4140 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1730889744
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1730889744
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1730889744
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1730889744
transform 1 0 6624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_74
timestamp 1730889744
transform 1 0 7912 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1730889744
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1730889744
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1730889744
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1730889744
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1730889744
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1730889744
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1730889744
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1730889744
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1730889744
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1730889744
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1730889744
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_35
timestamp 1730889744
transform 1 0 4324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1730889744
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_73
timestamp 1730889744
transform 1 0 7820 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1730889744
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_101
timestamp 1730889744
transform 1 0 10396 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_166
timestamp 1730889744
transform 1 0 16376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1730889744
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1730889744
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1730889744
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1730889744
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_205
timestamp 1730889744
transform 1 0 19964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1730889744
transform 1 0 20700 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_227
timestamp 1730889744
transform 1 0 21988 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1730889744
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1730889744
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_24
timestamp 1730889744
transform 1 0 3312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_30
timestamp 1730889744
transform 1 0 3864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_43
timestamp 1730889744
transform 1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1730889744
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1730889744
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1730889744
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1730889744
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1730889744
transform 1 0 13616 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1730889744
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1730889744
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1730889744
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_194
timestamp 1730889744
transform 1 0 18952 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_198
timestamp 1730889744
transform 1 0 19320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_216
timestamp 1730889744
transform 1 0 20976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_244
timestamp 1730889744
transform 1 0 23552 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_6
timestamp 1730889744
transform 1 0 1656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1730889744
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 1730889744
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_33
timestamp 1730889744
transform 1 0 4140 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1730889744
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_61
timestamp 1730889744
transform 1 0 6716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_69
timestamp 1730889744
transform 1 0 7452 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_76
timestamp 1730889744
transform 1 0 8096 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_101
timestamp 1730889744
transform 1 0 10396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_118
timestamp 1730889744
transform 1 0 11960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1730889744
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_168
timestamp 1730889744
transform 1 0 16560 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_178
timestamp 1730889744
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1730889744
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1730889744
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1730889744
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1730889744
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_217
timestamp 1730889744
transform 1 0 21068 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1730889744
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1730889744
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_9
timestamp 1730889744
transform 1 0 1932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_21
timestamp 1730889744
transform 1 0 3036 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_41
timestamp 1730889744
transform 1 0 4876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_47
timestamp 1730889744
transform 1 0 5428 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1730889744
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_65
timestamp 1730889744
transform 1 0 7084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_88
timestamp 1730889744
transform 1 0 9200 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1730889744
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1730889744
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_129
timestamp 1730889744
transform 1 0 12972 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1730889744
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1730889744
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1730889744
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_186
timestamp 1730889744
transform 1 0 18216 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1730889744
transform 1 0 18768 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_196
timestamp 1730889744
transform 1 0 19136 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_208
timestamp 1730889744
transform 1 0 20240 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_216
timestamp 1730889744
transform 1 0 20976 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1730889744
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_233
timestamp 1730889744
transform 1 0 22540 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1730889744
transform 1 0 23276 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1730889744
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1730889744
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1730889744
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1730889744
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1730889744
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1730889744
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_39
timestamp 1730889744
transform 1 0 4692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_64
timestamp 1730889744
transform 1 0 6992 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1730889744
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_92
timestamp 1730889744
transform 1 0 9568 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_100
timestamp 1730889744
transform 1 0 10304 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1730889744
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1730889744
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1730889744
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1730889744
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_234
timestamp 1730889744
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_246
timestamp 1730889744
transform 1 0 23736 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1730889744
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_30
timestamp 1730889744
transform 1 0 3864 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_44
timestamp 1730889744
transform 1 0 5152 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_95
timestamp 1730889744
transform 1 0 9844 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1730889744
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1730889744
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1730889744
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_199
timestamp 1730889744
transform 1 0 19412 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1730889744
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1730889744
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1730889744
transform 1 0 25760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1730889744
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1730889744
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1730889744
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1730889744
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_33
timestamp 1730889744
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_67
timestamp 1730889744
transform 1 0 7268 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_92
timestamp 1730889744
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_114
timestamp 1730889744
transform 1 0 11592 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1730889744
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_154
timestamp 1730889744
transform 1 0 15272 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_166
timestamp 1730889744
transform 1 0 16376 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1730889744
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_208
timestamp 1730889744
transform 1 0 20240 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_233
timestamp 1730889744
transform 1 0 22540 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1730889744
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1730889744
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_29
timestamp 1730889744
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_41
timestamp 1730889744
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1730889744
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1730889744
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_61
timestamp 1730889744
transform 1 0 6716 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_87
timestamp 1730889744
transform 1 0 9108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_95
timestamp 1730889744
transform 1 0 9844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_159
timestamp 1730889744
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1730889744
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1730889744
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1730889744
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_193
timestamp 1730889744
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_201
timestamp 1730889744
transform 1 0 19596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1730889744
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_238
timestamp 1730889744
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_242
timestamp 1730889744
transform 1 0 23368 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_3
timestamp 1730889744
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1730889744
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1730889744
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1730889744
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1730889744
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_58
timestamp 1730889744
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1730889744
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1730889744
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_97
timestamp 1730889744
transform 1 0 10028 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_128
timestamp 1730889744
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_149
timestamp 1730889744
transform 1 0 14812 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_161
timestamp 1730889744
transform 1 0 15916 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_168
timestamp 1730889744
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_181
timestamp 1730889744
transform 1 0 17756 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_185
timestamp 1730889744
transform 1 0 18124 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1730889744
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1730889744
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 1730889744
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_234
timestamp 1730889744
transform 1 0 22632 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1730889744
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1730889744
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_30
timestamp 1730889744
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1730889744
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_72
timestamp 1730889744
transform 1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_84
timestamp 1730889744
transform 1 0 8832 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_96
timestamp 1730889744
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_108
timestamp 1730889744
transform 1 0 11040 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_123
timestamp 1730889744
transform 1 0 12420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_151
timestamp 1730889744
transform 1 0 14996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1730889744
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1730889744
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_208
timestamp 1730889744
transform 1 0 20240 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1730889744
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1730889744
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1730889744
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_241
timestamp 1730889744
transform 1 0 23276 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1730889744
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_11
timestamp 1730889744
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1730889744
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1730889744
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_58
timestamp 1730889744
transform 1 0 6440 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1730889744
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1730889744
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_129
timestamp 1730889744
transform 1 0 12972 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1730889744
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_209
timestamp 1730889744
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_229
timestamp 1730889744
transform 1 0 22172 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp 1730889744
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1730889744
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_253
timestamp 1730889744
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1730889744
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_265
timestamp 1730889744
transform 1 0 25484 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1730889744
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1730889744
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1730889744
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_39
timestamp 1730889744
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1730889744
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1730889744
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1730889744
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1730889744
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp 1730889744
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_89
timestamp 1730889744
transform 1 0 9292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_145
timestamp 1730889744
transform 1 0 14444 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_149
timestamp 1730889744
transform 1 0 14812 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_157
timestamp 1730889744
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1730889744
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1730889744
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_211
timestamp 1730889744
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp 1730889744
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1730889744
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1730889744
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1730889744
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_261
timestamp 1730889744
transform 1 0 25116 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_269
timestamp 1730889744
transform 1 0 25852 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1730889744
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1730889744
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1730889744
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1730889744
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1730889744
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1730889744
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1730889744
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1730889744
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1730889744
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1730889744
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1730889744
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_103
timestamp 1730889744
transform 1 0 10580 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_112
timestamp 1730889744
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_146
timestamp 1730889744
transform 1 0 14536 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_158
timestamp 1730889744
transform 1 0 15640 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_164
timestamp 1730889744
transform 1 0 16192 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_168
timestamp 1730889744
transform 1 0 16560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1730889744
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1730889744
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_205
timestamp 1730889744
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_239
timestamp 1730889744
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1730889744
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1730889744
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1730889744
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_269
timestamp 1730889744
transform 1 0 25852 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1730889744
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1730889744
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1730889744
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1730889744
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1730889744
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1730889744
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1730889744
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1730889744
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1730889744
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1730889744
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_105
timestamp 1730889744
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1730889744
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_146
timestamp 1730889744
transform 1 0 14536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1730889744
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1730889744
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1730889744
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1730889744
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1730889744
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1730889744
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1730889744
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1730889744
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1730889744
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1730889744
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_261
timestamp 1730889744
transform 1 0 25116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 1730889744
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1730889744
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1730889744
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1730889744
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1730889744
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1730889744
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1730889744
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1730889744
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1730889744
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1730889744
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1730889744
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1730889744
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1730889744
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1730889744
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1730889744
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1730889744
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1730889744
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1730889744
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1730889744
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1730889744
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1730889744
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1730889744
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1730889744
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1730889744
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1730889744
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1730889744
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1730889744
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1730889744
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1730889744
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1730889744
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_269
timestamp 1730889744
transform 1 0 25852 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1730889744
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1730889744
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1730889744
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1730889744
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1730889744
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1730889744
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1730889744
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1730889744
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1730889744
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1730889744
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1730889744
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1730889744
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1730889744
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1730889744
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1730889744
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1730889744
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1730889744
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1730889744
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1730889744
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1730889744
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1730889744
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1730889744
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1730889744
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1730889744
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1730889744
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1730889744
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1730889744
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_261
timestamp 1730889744
transform 1 0 25116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_269
timestamp 1730889744
transform 1 0 25852 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1730889744
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1730889744
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1730889744
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1730889744
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1730889744
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1730889744
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1730889744
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1730889744
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1730889744
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1730889744
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1730889744
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1730889744
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1730889744
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1730889744
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1730889744
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1730889744
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1730889744
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1730889744
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1730889744
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1730889744
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1730889744
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1730889744
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1730889744
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1730889744
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1730889744
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1730889744
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1730889744
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1730889744
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1730889744
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1730889744
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1730889744
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1730889744
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_27
timestamp 1730889744
transform 1 0 3588 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_29
timestamp 1730889744
transform 1 0 3772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_41
timestamp 1730889744
transform 1 0 4876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1730889744
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1730889744
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1730889744
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_81
timestamp 1730889744
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_85
timestamp 1730889744
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_97
timestamp 1730889744
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1730889744
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1730889744
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1730889744
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_133
timestamp 1730889744
transform 1 0 13340 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_139
timestamp 1730889744
transform 1 0 13892 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_141
timestamp 1730889744
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_153
timestamp 1730889744
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1730889744
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1730889744
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1730889744
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_193
timestamp 1730889744
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_197
timestamp 1730889744
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_209
timestamp 1730889744
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1730889744
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1730889744
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1730889744
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_249
timestamp 1730889744
transform 1 0 24012 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1730889744
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1730889744
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_269
timestamp 1730889744
transform 1 0 25852 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 13248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1730889744
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1730889744
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1730889744
transform -1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1730889744
transform -1 0 25944 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1730889744
transform -1 0 25944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1730889744
transform -1 0 25944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1730889744
transform -1 0 25576 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1730889744
transform -1 0 25760 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1730889744
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1730889744
transform -1 0 12512 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1730889744
transform -1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1730889744
transform -1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1730889744
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1730889744
transform -1 0 25576 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1730889744
transform 1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1730889744
transform -1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1730889744
transform -1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1730889744
transform 1 0 12972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1730889744
transform -1 0 13432 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1730889744
transform -1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1730889744
transform 1 0 15824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1730889744
transform -1 0 18216 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1730889744
transform -1 0 13984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1730889744
transform -1 0 13616 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1730889744
transform -1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1730889744
transform -1 0 20700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1730889744
transform -1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1730889744
transform -1 0 20240 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1730889744
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1730889744
transform -1 0 18216 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1730889744
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1730889744
transform 1 0 15272 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1730889744
transform -1 0 19964 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1730889744
transform -1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1730889744
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1730889744
transform -1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1730889744
transform 1 0 11500 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1730889744
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1730889744
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1730889744
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1730889744
transform -1 0 16376 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1730889744
transform -1 0 12328 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1730889744
transform -1 0 18676 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1730889744
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1730889744
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1730889744
transform -1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1730889744
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1730889744
transform -1 0 18860 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1730889744
transform -1 0 13984 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1730889744
transform -1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1730889744
transform 1 0 19320 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1730889744
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1730889744
transform -1 0 14444 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1730889744
transform 1 0 18124 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1730889744
transform -1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1730889744
transform -1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1730889744
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1730889744
transform -1 0 25944 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1730889744
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1730889744
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 12328 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1730889744
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap66
timestamp 1730889744
transform 1 0 19964 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1730889744
transform 1 0 25576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1730889744
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1730889744
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1730889744
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1730889744
transform 1 0 25208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1730889744
transform 1 0 25576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1730889744
transform 1 0 25576 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1730889744
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1730889744
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1730889744
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1730889744
transform 1 0 25576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1730889744
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1730889744
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1730889744
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1730889744
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1730889744
transform 1 0 25208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1730889744
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1730889744
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1730889744
transform -1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1730889744
transform -1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1730889744
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1730889744
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1730889744
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1730889744
transform -1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1730889744
transform -1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1730889744
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1730889744
transform -1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1730889744
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1730889744
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1730889744
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1730889744
transform 1 0 25576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1730889744
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1730889744
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1730889744
transform 1 0 25576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1730889744
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1730889744
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1730889744
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1730889744
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1730889744
transform 1 0 25576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1730889744
transform 1 0 25576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1730889744
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1730889744
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1730889744
transform 1 0 25576 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1730889744
transform 1 0 25208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1730889744
transform -1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1730889744
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1730889744
transform -1 0 13984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1730889744
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1730889744
transform -1 0 16560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1730889744
transform -1 0 13340 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_46
timestamp 1730889744
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1730889744
transform -1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_47
timestamp 1730889744
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1730889744
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_48
timestamp 1730889744
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1730889744
transform -1 0 26220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_49
timestamp 1730889744
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1730889744
transform -1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_50
timestamp 1730889744
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1730889744
transform -1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_51
timestamp 1730889744
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1730889744
transform -1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_52
timestamp 1730889744
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1730889744
transform -1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_53
timestamp 1730889744
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1730889744
transform -1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_54
timestamp 1730889744
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1730889744
transform -1 0 26220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_55
timestamp 1730889744
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1730889744
transform -1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_56
timestamp 1730889744
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1730889744
transform -1 0 26220 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_57
timestamp 1730889744
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1730889744
transform -1 0 26220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_58
timestamp 1730889744
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1730889744
transform -1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_59
timestamp 1730889744
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1730889744
transform -1 0 26220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_60
timestamp 1730889744
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1730889744
transform -1 0 26220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_61
timestamp 1730889744
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1730889744
transform -1 0 26220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_62
timestamp 1730889744
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1730889744
transform -1 0 26220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_63
timestamp 1730889744
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1730889744
transform -1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_64
timestamp 1730889744
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1730889744
transform -1 0 26220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_65
timestamp 1730889744
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1730889744
transform -1 0 26220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_66
timestamp 1730889744
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1730889744
transform -1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_67
timestamp 1730889744
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1730889744
transform -1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_68
timestamp 1730889744
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1730889744
transform -1 0 26220 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_69
timestamp 1730889744
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1730889744
transform -1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_70
timestamp 1730889744
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1730889744
transform -1 0 26220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_71
timestamp 1730889744
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1730889744
transform -1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_72
timestamp 1730889744
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1730889744
transform -1 0 26220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_73
timestamp 1730889744
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1730889744
transform -1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_74
timestamp 1730889744
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1730889744
transform -1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_75
timestamp 1730889744
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1730889744
transform -1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_76
timestamp 1730889744
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1730889744
transform -1 0 26220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_77
timestamp 1730889744
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1730889744
transform -1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_78
timestamp 1730889744
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1730889744
transform -1 0 26220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_79
timestamp 1730889744
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1730889744
transform -1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_80
timestamp 1730889744
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1730889744
transform -1 0 26220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_81
timestamp 1730889744
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1730889744
transform -1 0 26220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_82
timestamp 1730889744
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1730889744
transform -1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_83
timestamp 1730889744
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1730889744
transform -1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_84
timestamp 1730889744
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1730889744
transform -1 0 26220 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_85
timestamp 1730889744
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1730889744
transform -1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_86
timestamp 1730889744
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1730889744
transform -1 0 26220 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_87
timestamp 1730889744
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1730889744
transform -1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_88
timestamp 1730889744
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1730889744
transform -1 0 26220 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_89
timestamp 1730889744
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1730889744
transform -1 0 26220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_90
timestamp 1730889744
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1730889744
transform -1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_91
timestamp 1730889744
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1730889744
transform -1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_92 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730889744
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_93
timestamp 1730889744
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp 1730889744
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp 1730889744
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp 1730889744
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_97
timestamp 1730889744
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 1730889744
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 1730889744
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1730889744
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_101
timestamp 1730889744
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_102
timestamp 1730889744
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_103
timestamp 1730889744
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_104
timestamp 1730889744
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_105
timestamp 1730889744
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_106
timestamp 1730889744
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_107
timestamp 1730889744
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_108
timestamp 1730889744
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_109
timestamp 1730889744
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_110
timestamp 1730889744
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_111
timestamp 1730889744
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_112
timestamp 1730889744
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_113
timestamp 1730889744
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_114
timestamp 1730889744
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_115
timestamp 1730889744
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_116
timestamp 1730889744
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_117
timestamp 1730889744
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_118
timestamp 1730889744
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_119
timestamp 1730889744
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_120
timestamp 1730889744
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_121
timestamp 1730889744
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_122
timestamp 1730889744
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_123
timestamp 1730889744
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_124
timestamp 1730889744
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_125
timestamp 1730889744
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_126
timestamp 1730889744
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_127
timestamp 1730889744
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_128
timestamp 1730889744
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_129
timestamp 1730889744
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_130
timestamp 1730889744
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_131
timestamp 1730889744
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1730889744
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_133
timestamp 1730889744
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_134
timestamp 1730889744
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_135
timestamp 1730889744
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_136
timestamp 1730889744
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1730889744
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_138
timestamp 1730889744
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_139
timestamp 1730889744
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_140
timestamp 1730889744
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1730889744
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1730889744
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1730889744
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_144
timestamp 1730889744
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_145
timestamp 1730889744
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1730889744
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1730889744
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1730889744
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_149
timestamp 1730889744
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1730889744
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1730889744
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1730889744
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1730889744
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1730889744
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1730889744
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1730889744
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1730889744
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1730889744
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_159
timestamp 1730889744
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1730889744
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1730889744
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1730889744
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1730889744
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_164
timestamp 1730889744
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_165
timestamp 1730889744
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1730889744
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1730889744
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_168
timestamp 1730889744
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_169
timestamp 1730889744
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_170
timestamp 1730889744
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1730889744
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1730889744
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_173
timestamp 1730889744
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_174
timestamp 1730889744
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_175
timestamp 1730889744
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_176
timestamp 1730889744
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1730889744
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_178
timestamp 1730889744
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_179
timestamp 1730889744
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_180
timestamp 1730889744
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_181
timestamp 1730889744
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 1730889744
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_183
timestamp 1730889744
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_184
timestamp 1730889744
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_185
timestamp 1730889744
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1730889744
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 1730889744
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 1730889744
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_189
timestamp 1730889744
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_190
timestamp 1730889744
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 1730889744
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 1730889744
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1730889744
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_194
timestamp 1730889744
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1730889744
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1730889744
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1730889744
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 1730889744
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 1730889744
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 1730889744
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 1730889744
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 1730889744
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 1730889744
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_204
timestamp 1730889744
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 1730889744
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1730889744
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1730889744
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 1730889744
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_209
timestamp 1730889744
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_210
timestamp 1730889744
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 1730889744
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 1730889744
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_213
timestamp 1730889744
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_214
timestamp 1730889744
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_215
timestamp 1730889744
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 1730889744
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 1730889744
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_218
timestamp 1730889744
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_219
timestamp 1730889744
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_220
timestamp 1730889744
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_221
timestamp 1730889744
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_222
timestamp 1730889744
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_223
timestamp 1730889744
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_224
timestamp 1730889744
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_225
timestamp 1730889744
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_226
timestamp 1730889744
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_227
timestamp 1730889744
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_228
timestamp 1730889744
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_229
timestamp 1730889744
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_230
timestamp 1730889744
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_231
timestamp 1730889744
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_232
timestamp 1730889744
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_233
timestamp 1730889744
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_234
timestamp 1730889744
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_235
timestamp 1730889744
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_236
timestamp 1730889744
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_237
timestamp 1730889744
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_238
timestamp 1730889744
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_239
timestamp 1730889744
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_240
timestamp 1730889744
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_241
timestamp 1730889744
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_242
timestamp 1730889744
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_243
timestamp 1730889744
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_244
timestamp 1730889744
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_245
timestamp 1730889744
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_246
timestamp 1730889744
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_247
timestamp 1730889744
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_248
timestamp 1730889744
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_249
timestamp 1730889744
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_250
timestamp 1730889744
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_251
timestamp 1730889744
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_252
timestamp 1730889744
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_253
timestamp 1730889744
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_254
timestamp 1730889744
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_255
timestamp 1730889744
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_256
timestamp 1730889744
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_257
timestamp 1730889744
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_258
timestamp 1730889744
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_259
timestamp 1730889744
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_260
timestamp 1730889744
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_261
timestamp 1730889744
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_262
timestamp 1730889744
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_263
timestamp 1730889744
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_264
timestamp 1730889744
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_265
timestamp 1730889744
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_266
timestamp 1730889744
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_267
timestamp 1730889744
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_268
timestamp 1730889744
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_269
timestamp 1730889744
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_270
timestamp 1730889744
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_271
timestamp 1730889744
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_272
timestamp 1730889744
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_273
timestamp 1730889744
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_274
timestamp 1730889744
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_275
timestamp 1730889744
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_276
timestamp 1730889744
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_277
timestamp 1730889744
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_278
timestamp 1730889744
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_279
timestamp 1730889744
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_280
timestamp 1730889744
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_281
timestamp 1730889744
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_282
timestamp 1730889744
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_283
timestamp 1730889744
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_284
timestamp 1730889744
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_285
timestamp 1730889744
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_286
timestamp 1730889744
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_287
timestamp 1730889744
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_288
timestamp 1730889744
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_289
timestamp 1730889744
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_290
timestamp 1730889744
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_291
timestamp 1730889744
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_292
timestamp 1730889744
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_293
timestamp 1730889744
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_294
timestamp 1730889744
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_295
timestamp 1730889744
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_296
timestamp 1730889744
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_297
timestamp 1730889744
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_298
timestamp 1730889744
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_299
timestamp 1730889744
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_300
timestamp 1730889744
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_301
timestamp 1730889744
transform 1 0 8832 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_302
timestamp 1730889744
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_303
timestamp 1730889744
transform 1 0 13984 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_304
timestamp 1730889744
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_305
timestamp 1730889744
transform 1 0 19136 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_306
timestamp 1730889744
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_307
timestamp 1730889744
transform 1 0 24288 0 -1 27200
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 27248 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 27248 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 b0
port 2 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 b1
port 3 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 clk
port 4 nsew signal input
flabel metal3 s 26532 22448 27332 22568 0 FreeSans 480 0 0 0 compr
port 5 nsew signal input
flabel metal3 s 26532 21768 27332 21888 0 FreeSans 480 0 0 0 dac[0]
port 6 nsew signal output
flabel metal3 s 26532 21088 27332 21208 0 FreeSans 480 0 0 0 dac[1]
port 7 nsew signal output
flabel metal3 s 26532 19728 27332 19848 0 FreeSans 480 0 0 0 dac[2]
port 8 nsew signal output
flabel metal3 s 26532 17008 27332 17128 0 FreeSans 480 0 0 0 dac[3]
port 9 nsew signal output
flabel metal3 s 26532 19048 27332 19168 0 FreeSans 480 0 0 0 dac[4]
port 10 nsew signal output
flabel metal3 s 26532 17688 27332 17808 0 FreeSans 480 0 0 0 dac[5]
port 11 nsew signal output
flabel metal3 s 26532 20408 27332 20528 0 FreeSans 480 0 0 0 dac[6]
port 12 nsew signal output
flabel metal3 s 26532 14968 27332 15088 0 FreeSans 480 0 0 0 dac[7]
port 13 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dac_coupl
port 14 nsew signal output
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 m0
port 15 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 m1
port 16 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 reg0[0]
port 17 nsew signal output
flabel metal3 s 26532 12928 27332 13048 0 FreeSans 480 0 0 0 reg0[1]
port 18 nsew signal output
flabel metal3 s 26532 2728 27332 2848 0 FreeSans 480 0 0 0 reg0[2]
port 19 nsew signal output
flabel metal3 s 26532 3408 27332 3528 0 FreeSans 480 0 0 0 reg0[3]
port 20 nsew signal output
flabel metal3 s 26532 15648 27332 15768 0 FreeSans 480 0 0 0 reg0[4]
port 21 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 reg0[5]
port 22 nsew signal output
flabel metal3 s 26532 4088 27332 4208 0 FreeSans 480 0 0 0 reg0[6]
port 23 nsew signal output
flabel metal3 s 26532 6808 27332 6928 0 FreeSans 480 0 0 0 reg0[7]
port 24 nsew signal output
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 reg1[0]
port 25 nsew signal output
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 reg1[1]
port 26 nsew signal output
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 reg1[2]
port 27 nsew signal output
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 reg1[3]
port 28 nsew signal output
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 reg1[4]
port 29 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 reg1[5]
port 30 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 reg1[6]
port 31 nsew signal output
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 reg1[7]
port 32 nsew signal output
flabel metal3 s 26532 4768 27332 4888 0 FreeSans 480 0 0 0 reg2[0]
port 33 nsew signal output
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 reg2[1]
port 34 nsew signal output
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 reg2[2]
port 35 nsew signal output
flabel metal3 s 26532 5448 27332 5568 0 FreeSans 480 0 0 0 reg2[3]
port 36 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 reg2[4]
port 37 nsew signal output
flabel metal3 s 26532 6128 27332 6248 0 FreeSans 480 0 0 0 reg2[5]
port 38 nsew signal output
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 reg2[6]
port 39 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 reg2[7]
port 40 nsew signal output
flabel metal3 s 26532 8848 27332 8968 0 FreeSans 480 0 0 0 reg3[0]
port 41 nsew signal output
flabel metal3 s 26532 10208 27332 10328 0 FreeSans 480 0 0 0 reg3[1]
port 42 nsew signal output
flabel metal3 s 26532 10888 27332 11008 0 FreeSans 480 0 0 0 reg3[2]
port 43 nsew signal output
flabel metal3 s 26532 7488 27332 7608 0 FreeSans 480 0 0 0 reg3[3]
port 44 nsew signal output
flabel metal3 s 26532 12248 27332 12368 0 FreeSans 480 0 0 0 reg3[4]
port 45 nsew signal output
flabel metal3 s 26532 8168 27332 8288 0 FreeSans 480 0 0 0 reg3[5]
port 46 nsew signal output
flabel metal3 s 26532 11568 27332 11688 0 FreeSans 480 0 0 0 reg3[6]
port 47 nsew signal output
flabel metal3 s 26532 9528 27332 9648 0 FreeSans 480 0 0 0 reg3[7]
port 48 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 reg4[0]
port 49 nsew signal output
flabel metal3 s 26532 14288 27332 14408 0 FreeSans 480 0 0 0 reg4[1]
port 50 nsew signal output
flabel metal3 s 26532 13608 27332 13728 0 FreeSans 480 0 0 0 reg4[2]
port 51 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 reg4[3]
port 52 nsew signal output
flabel metal3 s 26532 16328 27332 16448 0 FreeSans 480 0 0 0 reg4[4]
port 53 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 reg4[5]
port 54 nsew signal output
flabel metal3 s 26532 18368 27332 18488 0 FreeSans 480 0 0 0 reg4[6]
port 55 nsew signal output
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 reg4[7]
port 56 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 rst
port 57 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 rx
port 58 nsew signal input
flabel metal2 s 12898 28676 12954 29476 0 FreeSans 224 90 0 0 tx
port 59 nsew signal output
rlabel metal1 13662 27200 13662 27200 0 VGND
rlabel metal1 13662 26656 13662 26656 0 VPWR
rlabel metal2 15410 10914 15410 10914 0 _0000_
rlabel metal2 24702 20706 24702 20706 0 _0001_
rlabel metal1 1927 17578 1927 17578 0 _0002_
rlabel via1 2994 18258 2994 18258 0 _0003_
rlabel metal1 2116 20570 2116 20570 0 _0004_
rlabel metal2 2162 21726 2162 21726 0 _0005_
rlabel metal2 2530 22882 2530 22882 0 _0006_
rlabel viali 4917 22610 4917 22610 0 _0007_
rlabel metal1 5423 23086 5423 23086 0 _0008_
rlabel metal2 7038 22882 7038 22882 0 _0009_
rlabel metal2 8234 21692 8234 21692 0 _0010_
rlabel metal2 8418 20434 8418 20434 0 _0011_
rlabel metal1 10038 18258 10038 18258 0 _0012_
rlabel via1 10078 17646 10078 17646 0 _0013_
rlabel metal1 9200 17850 9200 17850 0 _0014_
rlabel via1 10805 5678 10805 5678 0 _0015_
rlabel metal1 12834 13804 12834 13804 0 _0016_
rlabel metal1 13519 4114 13519 4114 0 _0017_
rlabel metal2 21206 13090 21206 13090 0 _0018_
rlabel metal1 19964 11322 19964 11322 0 _0019_
rlabel metal1 13059 4590 13059 4590 0 _0020_
rlabel metal2 21390 14144 21390 14144 0 _0021_
rlabel metal2 14122 6086 14122 6086 0 _0022_
rlabel metal1 20286 13498 20286 13498 0 _0023_
rlabel metal1 15502 6426 15502 6426 0 _0024_
rlabel metal1 24042 8534 24042 8534 0 _0025_
rlabel metal1 24242 11152 24242 11152 0 _0026_
rlabel metal1 24226 10710 24226 10710 0 _0027_
rlabel metal1 24042 7446 24042 7446 0 _0028_
rlabel metal1 24697 12818 24697 12818 0 _0029_
rlabel metal1 23966 7310 23966 7310 0 _0030_
rlabel metal1 21850 11322 21850 11322 0 _0031_
rlabel metal1 20868 8874 20868 8874 0 _0032_
rlabel metal1 24456 4522 24456 4522 0 _0033_
rlabel metal1 24932 3706 24932 3706 0 _0034_
rlabel via1 22949 3094 22949 3094 0 _0035_
rlabel metal1 24318 5270 24318 5270 0 _0036_
rlabel via1 22489 3502 22489 3502 0 _0037_
rlabel metal1 23766 6358 23766 6358 0 _0038_
rlabel metal2 21850 3298 21850 3298 0 _0039_
rlabel metal1 21942 5168 21942 5168 0 _0040_
rlabel via1 14393 3434 14393 3434 0 _0041_
rlabel metal1 17705 3434 17705 3434 0 _0042_
rlabel metal2 19274 3910 19274 3910 0 _0043_
rlabel metal1 14577 3094 14577 3094 0 _0044_
rlabel metal1 19197 3094 19197 3094 0 _0045_
rlabel metal1 15824 5338 15824 5338 0 _0046_
rlabel metal2 16698 3298 16698 3298 0 _0047_
rlabel metal2 18078 4998 18078 4998 0 _0048_
rlabel metal1 19304 6698 19304 6698 0 _0049_
rlabel metal1 24456 13226 24456 13226 0 _0050_
rlabel metal1 23950 9622 23950 9622 0 _0051_
rlabel metal1 21201 5610 21201 5610 0 _0052_
rlabel metal2 24334 14178 24334 14178 0 _0053_
rlabel via1 19361 6358 19361 6358 0 _0054_
rlabel metal1 21104 10030 21104 10030 0 _0055_
rlabel metal1 20930 7514 20930 7514 0 _0056_
rlabel metal1 15419 14314 15419 14314 0 _0057_
rlabel metal2 17894 13090 17894 13090 0 _0058_
rlabel metal1 18073 11118 18073 11118 0 _0059_
rlabel metal1 15502 13498 15502 13498 0 _0060_
rlabel metal2 18630 14178 18630 14178 0 _0061_
rlabel metal1 13984 13498 13984 13498 0 _0062_
rlabel metal1 18441 13974 18441 13974 0 _0063_
rlabel metal1 16371 14314 16371 14314 0 _0064_
rlabel via1 17889 10030 17889 10030 0 _0065_
rlabel metal1 18579 9622 18579 9622 0 _0066_
rlabel via1 17337 11798 17337 11798 0 _0067_
rlabel metal1 15359 9622 15359 9622 0 _0068_
rlabel metal1 16003 8942 16003 8942 0 _0069_
rlabel metal2 8786 22746 8786 22746 0 _0070_
rlabel metal2 10534 23494 10534 23494 0 _0071_
rlabel metal1 12190 23222 12190 23222 0 _0072_
rlabel metal1 11454 23154 11454 23154 0 _0073_
rlabel metal1 12634 24106 12634 24106 0 _0074_
rlabel metal2 14858 19618 14858 19618 0 _0075_
rlabel metal2 11822 16966 11822 16966 0 _0076_
rlabel metal2 12098 15878 12098 15878 0 _0077_
rlabel metal1 12742 15912 12742 15912 0 _0078_
rlabel metal1 15425 17578 15425 17578 0 _0079_
rlabel metal1 15328 17170 15328 17170 0 _0080_
rlabel via1 15598 18326 15598 18326 0 _0081_
rlabel metal1 14904 21114 14904 21114 0 _0082_
rlabel metal1 2336 4590 2336 4590 0 _0083_
rlabel metal1 4012 5202 4012 5202 0 _0084_
rlabel metal2 2346 6562 2346 6562 0 _0085_
rlabel via1 2341 7378 2341 7378 0 _0086_
rlabel via1 2810 8942 2810 8942 0 _0087_
rlabel viali 3169 8466 3169 8466 0 _0088_
rlabel metal2 5658 8262 5658 8262 0 _0089_
rlabel metal1 7318 5678 7318 5678 0 _0090_
rlabel metal2 5566 5474 5566 5474 0 _0091_
rlabel metal1 8882 5202 8882 5202 0 _0092_
rlabel metal1 9802 5610 9802 5610 0 _0093_
rlabel metal1 8142 6222 8142 6222 0 _0094_
rlabel via1 10253 9554 10253 9554 0 _0095_
rlabel metal1 8408 8466 8408 8466 0 _0096_
rlabel metal1 9506 8874 9506 8874 0 _0097_
rlabel metal1 10411 7786 10411 7786 0 _0098_
rlabel metal1 11392 19414 11392 19414 0 _0099_
rlabel via1 12654 20502 12654 20502 0 _0100_
rlabel metal1 12972 20570 12972 20570 0 _0101_
rlabel via1 10161 20910 10161 20910 0 _0102_
rlabel metal1 10897 21522 10897 21522 0 _0103_
rlabel via1 1881 13906 1881 13906 0 _0104_
rlabel metal1 3158 15062 3158 15062 0 _0105_
rlabel metal2 2438 15878 2438 15878 0 _0106_
rlabel metal2 2162 13906 2162 13906 0 _0107_
rlabel via1 1973 11730 1973 11730 0 _0108_
rlabel metal2 3266 11560 3266 11560 0 _0109_
rlabel metal1 4104 10642 4104 10642 0 _0110_
rlabel metal1 5612 10778 5612 10778 0 _0111_
rlabel metal1 8606 10710 8606 10710 0 _0112_
rlabel metal1 8832 11322 8832 11322 0 _0113_
rlabel metal1 9756 12886 9756 12886 0 _0114_
rlabel metal1 9046 14314 9046 14314 0 _0115_
rlabel metal1 9292 13702 9292 13702 0 _0116_
rlabel via1 24053 17170 24053 17170 0 _0117_
rlabel metal1 12673 12342 12673 12342 0 _0118_
rlabel metal1 18001 20502 18001 20502 0 _0119_
rlabel metal1 19335 19754 19335 19754 0 _0120_
rlabel metal1 18119 16150 18119 16150 0 _0121_
rlabel metal1 18185 18326 18185 18326 0 _0122_
rlabel via1 19738 16082 19738 16082 0 _0123_
rlabel metal1 21492 16082 21492 16082 0 _0124_
rlabel metal1 17981 16558 17981 16558 0 _0125_
rlabel metal2 24426 22406 24426 22406 0 _0126_
rlabel metal1 24150 21114 24150 21114 0 _0127_
rlabel metal1 24283 19414 24283 19414 0 _0128_
rlabel metal1 24456 16490 24456 16490 0 _0129_
rlabel metal2 23322 15266 23322 15266 0 _0130_
rlabel metal1 21436 23834 21436 23834 0 _0131_
rlabel metal2 21114 23698 21114 23698 0 _0132_
rlabel metal1 19228 23290 19228 23290 0 _0133_
rlabel metal1 12001 9622 12001 9622 0 _0134_
rlabel metal2 12926 12070 12926 12070 0 _0135_
rlabel metal1 11914 11322 11914 11322 0 _0136_
rlabel metal1 16325 19822 16325 19822 0 _0137_
rlabel metal1 16008 22746 16008 22746 0 _0138_
rlabel via1 14117 8466 14117 8466 0 _0139_
rlabel metal1 15313 11730 15313 11730 0 _0140_
rlabel metal1 16688 23086 16688 23086 0 _0141_
rlabel metal1 18308 24378 18308 24378 0 _0142_
rlabel metal1 14152 7786 14152 7786 0 _0143_
rlabel metal1 14628 11866 14628 11866 0 _0144_
rlabel metal1 18124 22746 18124 22746 0 _0145_
rlabel metal1 24237 18326 24237 18326 0 _0146_
rlabel metal2 10902 24174 10902 24174 0 _0147_
rlabel metal2 20194 16864 20194 16864 0 _0148_
rlabel metal2 18722 8704 18722 8704 0 _0149_
rlabel metal2 19090 8636 19090 8636 0 _0150_
rlabel metal2 17894 23222 17894 23222 0 _0151_
rlabel metal2 18998 22406 18998 22406 0 _0152_
rlabel metal1 21574 21352 21574 21352 0 _0153_
rlabel metal1 6992 13294 6992 13294 0 _0154_
rlabel metal2 8142 6528 8142 6528 0 _0155_
rlabel metal1 20792 15674 20792 15674 0 _0156_
rlabel metal2 3634 14926 3634 14926 0 _0157_
rlabel via2 11638 7259 11638 7259 0 _0158_
rlabel metal1 13294 8908 13294 8908 0 _0159_
rlabel metal2 12466 9724 12466 9724 0 _0160_
rlabel metal2 13202 10948 13202 10948 0 _0161_
rlabel metal1 13432 7922 13432 7922 0 _0162_
rlabel metal1 10718 7242 10718 7242 0 _0163_
rlabel metal1 11914 10506 11914 10506 0 _0164_
rlabel metal2 6578 15674 6578 15674 0 _0165_
rlabel metal1 7991 13362 7991 13362 0 _0166_
rlabel metal1 8050 13294 8050 13294 0 _0167_
rlabel metal2 7866 13498 7866 13498 0 _0168_
rlabel metal1 5980 8806 5980 8806 0 _0169_
rlabel metal1 7498 17102 7498 17102 0 _0170_
rlabel metal1 7636 13294 7636 13294 0 _0171_
rlabel metal1 7452 13906 7452 13906 0 _0172_
rlabel metal1 5980 16218 5980 16218 0 _0173_
rlabel metal1 4600 19278 4600 19278 0 _0174_
rlabel metal2 5842 20978 5842 20978 0 _0175_
rlabel metal2 3910 19550 3910 19550 0 _0176_
rlabel metal1 5796 13294 5796 13294 0 _0177_
rlabel metal1 5198 11866 5198 11866 0 _0178_
rlabel metal1 6118 13328 6118 13328 0 _0179_
rlabel metal1 6072 13974 6072 13974 0 _0180_
rlabel metal1 4922 14416 4922 14416 0 _0181_
rlabel metal1 5198 13294 5198 13294 0 _0182_
rlabel metal2 4738 15130 4738 15130 0 _0183_
rlabel metal2 5842 14110 5842 14110 0 _0184_
rlabel metal1 5428 15062 5428 15062 0 _0185_
rlabel metal1 5290 15028 5290 15028 0 _0186_
rlabel metal2 6118 14620 6118 14620 0 _0187_
rlabel metal1 5934 13872 5934 13872 0 _0188_
rlabel metal1 5658 12682 5658 12682 0 _0189_
rlabel metal2 5474 13838 5474 13838 0 _0190_
rlabel metal1 5888 13430 5888 13430 0 _0191_
rlabel metal1 5244 13498 5244 13498 0 _0192_
rlabel metal1 6118 13804 6118 13804 0 _0193_
rlabel metal1 8418 13362 8418 13362 0 _0194_
rlabel metal1 8142 13498 8142 13498 0 _0195_
rlabel metal2 8050 14178 8050 14178 0 _0196_
rlabel metal1 10258 15504 10258 15504 0 _0197_
rlabel metal1 6486 14382 6486 14382 0 _0198_
rlabel metal1 6540 13974 6540 13974 0 _0199_
rlabel metal1 6946 13906 6946 13906 0 _0200_
rlabel metal1 8142 12614 8142 12614 0 _0201_
rlabel metal1 14306 10608 14306 10608 0 _0202_
rlabel metal1 14674 10778 14674 10778 0 _0203_
rlabel metal2 15962 10778 15962 10778 0 _0204_
rlabel metal2 15548 19108 15548 19108 0 _0205_
rlabel metal1 19550 20876 19550 20876 0 _0206_
rlabel metal1 16192 21998 16192 21998 0 _0207_
rlabel metal1 21298 21590 21298 21590 0 _0208_
rlabel viali 21114 20911 21114 20911 0 _0209_
rlabel metal1 20838 21454 20838 21454 0 _0210_
rlabel metal1 21620 22746 21620 22746 0 _0211_
rlabel metal1 21436 18734 21436 18734 0 _0212_
rlabel metal2 21850 16762 21850 16762 0 _0213_
rlabel metal1 22310 21862 22310 21862 0 _0214_
rlabel metal2 23598 16524 23598 16524 0 _0215_
rlabel metal1 21482 19448 21482 19448 0 _0216_
rlabel via1 12466 13685 12466 13685 0 _0217_
rlabel metal2 12006 7072 12006 7072 0 _0218_
rlabel metal2 17342 14722 17342 14722 0 _0219_
rlabel metal1 19918 21522 19918 21522 0 _0220_
rlabel metal1 21896 19346 21896 19346 0 _0221_
rlabel metal1 22034 20400 22034 20400 0 _0222_
rlabel metal2 20010 21250 20010 21250 0 _0223_
rlabel metal1 19504 20774 19504 20774 0 _0224_
rlabel metal2 21390 20825 21390 20825 0 _0225_
rlabel metal1 23598 20366 23598 20366 0 _0226_
rlabel metal1 23000 20910 23000 20910 0 _0227_
rlabel metal1 23736 20298 23736 20298 0 _0228_
rlabel metal2 7682 17238 7682 17238 0 _0229_
rlabel metal2 7590 17884 7590 17884 0 _0230_
rlabel metal1 7314 17272 7314 17272 0 _0231_
rlabel metal2 5842 18445 5842 18445 0 _0232_
rlabel metal1 4508 18326 4508 18326 0 _0233_
rlabel metal2 4462 18428 4462 18428 0 _0234_
rlabel metal2 5106 18836 5106 18836 0 _0235_
rlabel metal1 5612 19822 5612 19822 0 _0236_
rlabel metal1 5934 19822 5934 19822 0 _0237_
rlabel metal1 6624 20026 6624 20026 0 _0238_
rlabel metal1 5842 19346 5842 19346 0 _0239_
rlabel metal1 5152 19142 5152 19142 0 _0240_
rlabel metal2 4738 19040 4738 19040 0 _0241_
rlabel metal2 6026 18700 6026 18700 0 _0242_
rlabel via1 6923 19346 6923 19346 0 _0243_
rlabel metal1 5382 19856 5382 19856 0 _0244_
rlabel metal2 4646 20604 4646 20604 0 _0245_
rlabel metal2 5658 19244 5658 19244 0 _0246_
rlabel metal2 5198 20026 5198 20026 0 _0247_
rlabel metal1 5566 18598 5566 18598 0 _0248_
rlabel viali 6486 19346 6486 19346 0 _0249_
rlabel metal1 6900 18190 6900 18190 0 _0250_
rlabel metal1 6808 17782 6808 17782 0 _0251_
rlabel metal1 5658 17680 5658 17680 0 _0252_
rlabel metal1 7222 17850 7222 17850 0 _0253_
rlabel metal1 8648 19414 8648 19414 0 _0254_
rlabel metal1 5428 17850 5428 17850 0 _0255_
rlabel metal2 5934 18428 5934 18428 0 _0256_
rlabel metal1 8234 18394 8234 18394 0 _0257_
rlabel metal2 2622 18972 2622 18972 0 _0258_
rlabel metal1 1794 20366 1794 20366 0 _0259_
rlabel metal2 1978 20230 1978 20230 0 _0260_
rlabel metal1 2057 20366 2057 20366 0 _0261_
rlabel metal1 5428 21998 5428 21998 0 _0262_
rlabel metal2 3358 21318 3358 21318 0 _0263_
rlabel metal2 3634 21794 3634 21794 0 _0264_
rlabel metal1 3266 22576 3266 22576 0 _0265_
rlabel metal1 4692 21998 4692 21998 0 _0266_
rlabel metal1 4830 21930 4830 21930 0 _0267_
rlabel metal1 4784 22202 4784 22202 0 _0268_
rlabel metal1 6854 21488 6854 21488 0 _0269_
rlabel metal1 6118 22032 6118 22032 0 _0270_
rlabel metal1 5716 23630 5716 23630 0 _0271_
rlabel metal1 7071 22542 7071 22542 0 _0272_
rlabel metal1 8832 21998 8832 21998 0 _0273_
rlabel metal2 7130 21692 7130 21692 0 _0274_
rlabel metal1 8246 21930 8246 21930 0 _0275_
rlabel metal1 8510 19856 8510 19856 0 _0276_
rlabel metal2 8694 20026 8694 20026 0 _0277_
rlabel metal1 8430 19754 8430 19754 0 _0278_
rlabel metal1 8556 17102 8556 17102 0 _0279_
rlabel via1 10337 18326 10337 18326 0 _0280_
rlabel metal1 8464 17306 8464 17306 0 _0281_
rlabel metal1 8660 17714 8660 17714 0 _0282_
rlabel metal2 11362 6426 11362 6426 0 _0283_
rlabel metal2 13110 14450 13110 14450 0 _0284_
rlabel metal1 12850 13974 12850 13974 0 _0285_
rlabel metal1 17710 7752 17710 7752 0 _0286_
rlabel metal2 21298 7378 21298 7378 0 _0287_
rlabel metal2 21850 13770 21850 13770 0 _0288_
rlabel metal2 20562 13345 20562 13345 0 _0289_
rlabel metal2 14582 5066 14582 5066 0 _0290_
rlabel metal1 20746 12852 20746 12852 0 _0291_
rlabel metal2 20470 11594 20470 11594 0 _0292_
rlabel metal1 13754 5236 13754 5236 0 _0293_
rlabel metal1 20930 14416 20930 14416 0 _0294_
rlabel metal2 14582 6154 14582 6154 0 _0295_
rlabel metal2 21298 13056 21298 13056 0 _0296_
rlabel metal2 16054 6460 16054 6460 0 _0297_
rlabel metal1 22908 12410 22908 12410 0 _0298_
rlabel metal1 22908 11050 22908 11050 0 _0299_
rlabel metal1 23690 10710 23690 10710 0 _0300_
rlabel metal1 23322 8432 23322 8432 0 _0301_
rlabel metal1 23782 11084 23782 11084 0 _0302_
rlabel metal2 23598 10948 23598 10948 0 _0303_
rlabel metal1 23414 7820 23414 7820 0 _0304_
rlabel metal1 24610 12172 24610 12172 0 _0305_
rlabel metal2 23506 7038 23506 7038 0 _0306_
rlabel metal1 22218 11152 22218 11152 0 _0307_
rlabel metal1 20838 9044 20838 9044 0 _0308_
rlabel metal2 20286 7140 20286 7140 0 _0309_
rlabel metal1 21160 2414 21160 2414 0 _0310_
rlabel metal1 21390 5236 21390 5236 0 _0311_
rlabel metal2 23782 5202 23782 5202 0 _0312_
rlabel metal2 24518 3332 24518 3332 0 _0313_
rlabel metal1 23644 3706 23644 3706 0 _0314_
rlabel metal1 23552 5202 23552 5202 0 _0315_
rlabel metal1 21988 4114 21988 4114 0 _0316_
rlabel metal1 23506 5882 23506 5882 0 _0317_
rlabel metal1 21942 2550 21942 2550 0 _0318_
rlabel metal1 21574 4794 21574 4794 0 _0319_
rlabel metal2 18262 5474 18262 5474 0 _0320_
rlabel metal1 18722 2482 18722 2482 0 _0321_
rlabel metal1 20010 4080 20010 4080 0 _0322_
rlabel metal1 15502 3094 15502 3094 0 _0323_
rlabel metal1 17434 3162 17434 3162 0 _0324_
rlabel metal2 19826 3315 19826 3315 0 _0325_
rlabel metal1 15410 3162 15410 3162 0 _0326_
rlabel metal1 19458 2346 19458 2346 0 _0327_
rlabel metal1 16238 5236 16238 5236 0 _0328_
rlabel metal1 17158 3094 17158 3094 0 _0329_
rlabel metal1 18538 4556 18538 4556 0 _0330_
rlabel metal2 16238 4318 16238 4318 0 _0331_
rlabel metal1 20378 7310 20378 7310 0 _0332_
rlabel metal1 21390 10608 21390 10608 0 _0333_
rlabel metal2 18630 6834 18630 6834 0 _0334_
rlabel metal1 23782 13328 23782 13328 0 _0335_
rlabel metal1 24058 9146 24058 9146 0 _0336_
rlabel metal2 20930 6970 20930 6970 0 _0337_
rlabel metal1 23874 13872 23874 13872 0 _0338_
rlabel metal1 19366 7412 19366 7412 0 _0339_
rlabel metal1 21482 10676 21482 10676 0 _0340_
rlabel metal1 21298 7344 21298 7344 0 _0341_
rlabel metal1 15686 4794 15686 4794 0 _0342_
rlabel metal1 20102 5032 20102 5032 0 _0343_
rlabel metal1 15732 15062 15732 15062 0 _0344_
rlabel metal1 20470 3366 20470 3366 0 _0345_
rlabel metal1 20608 12342 20608 12342 0 _0346_
rlabel metal1 18998 12818 18998 12818 0 _0347_
rlabel metal1 21068 3910 21068 3910 0 _0348_
rlabel metal1 23000 10234 23000 10234 0 _0349_
rlabel metal2 18998 11458 18998 11458 0 _0350_
rlabel metal2 15410 5729 15410 5729 0 _0351_
rlabel metal1 15778 3978 15778 3978 0 _0352_
rlabel metal1 15226 13226 15226 13226 0 _0353_
rlabel metal1 20654 12784 20654 12784 0 _0354_
rlabel metal1 19826 12750 19826 12750 0 _0355_
rlabel metal2 19550 13430 19550 13430 0 _0356_
rlabel metal1 16330 6426 16330 6426 0 _0357_
rlabel metal1 18814 6392 18814 6392 0 _0358_
rlabel metal1 13892 13226 13892 13226 0 _0359_
rlabel metal1 21022 12240 21022 12240 0 _0360_
rlabel metal1 21298 3162 21298 3162 0 _0361_
rlabel metal1 20056 13906 20056 13906 0 _0362_
rlabel metal2 20010 6120 20010 6120 0 _0363_
rlabel metal1 17250 7344 17250 7344 0 _0364_
rlabel metal1 16974 14926 16974 14926 0 _0365_
rlabel metal1 15962 10132 15962 10132 0 _0366_
rlabel metal1 17250 9554 17250 9554 0 _0367_
rlabel metal1 11546 23290 11546 23290 0 _0368_
rlabel metal1 12604 23086 12604 23086 0 _0369_
rlabel metal1 13294 23120 13294 23120 0 _0370_
rlabel metal1 13708 22950 13708 22950 0 _0371_
rlabel metal1 12006 24038 12006 24038 0 _0372_
rlabel metal1 13524 21114 13524 21114 0 _0373_
rlabel metal1 14076 23766 14076 23766 0 _0374_
rlabel via2 14030 20587 14030 20587 0 _0375_
rlabel metal2 11914 18326 11914 18326 0 _0376_
rlabel metal2 12650 18020 12650 18020 0 _0377_
rlabel metal1 12374 18258 12374 18258 0 _0378_
rlabel metal1 13018 18394 13018 18394 0 _0379_
rlabel metal1 13248 18258 13248 18258 0 _0380_
rlabel metal1 13478 18700 13478 18700 0 _0381_
rlabel metal2 13846 18666 13846 18666 0 _0382_
rlabel metal1 13294 17850 13294 17850 0 _0383_
rlabel metal1 13248 18734 13248 18734 0 _0384_
rlabel metal2 13018 18428 13018 18428 0 _0385_
rlabel metal1 13524 20230 13524 20230 0 _0386_
rlabel metal1 13708 18258 13708 18258 0 _0387_
rlabel via2 13570 18411 13570 18411 0 _0388_
rlabel metal1 12972 23086 12972 23086 0 _0389_
rlabel metal1 12558 21930 12558 21930 0 _0390_
rlabel metal2 16698 19142 16698 19142 0 _0391_
rlabel metal1 15134 15606 15134 15606 0 _0392_
rlabel metal1 13202 15402 13202 15402 0 _0393_
rlabel metal1 15824 15674 15824 15674 0 _0394_
rlabel metal1 16100 16762 16100 16762 0 _0395_
rlabel metal1 16928 17034 16928 17034 0 _0396_
rlabel metal2 17894 18258 17894 18258 0 _0397_
rlabel metal2 15226 20672 15226 20672 0 _0398_
rlabel metal1 5658 7854 5658 7854 0 _0399_
rlabel metal2 4646 5168 4646 5168 0 _0400_
rlabel metal1 4002 6426 4002 6426 0 _0401_
rlabel metal2 4370 7650 4370 7650 0 _0402_
rlabel metal1 4784 7922 4784 7922 0 _0403_
rlabel metal1 4784 7854 4784 7854 0 _0404_
rlabel metal1 5014 7820 5014 7820 0 _0405_
rlabel metal1 6982 7378 6982 7378 0 _0406_
rlabel metal2 9154 7650 9154 7650 0 _0407_
rlabel metal2 7130 7548 7130 7548 0 _0408_
rlabel metal1 7268 7378 7268 7378 0 _0409_
rlabel metal1 7452 7378 7452 7378 0 _0410_
rlabel metal1 7544 8058 7544 8058 0 _0411_
rlabel metal1 7866 7718 7866 7718 0 _0412_
rlabel metal2 5842 6528 5842 6528 0 _0413_
rlabel metal1 3851 5338 3851 5338 0 _0414_
rlabel metal1 2254 6392 2254 6392 0 _0415_
rlabel metal2 3634 8466 3634 8466 0 _0416_
rlabel metal2 2806 7242 2806 7242 0 _0417_
rlabel metal1 3174 7990 3174 7990 0 _0418_
rlabel metal2 1794 9112 1794 9112 0 _0419_
rlabel metal1 4140 8466 4140 8466 0 _0420_
rlabel metal2 3174 8160 3174 8160 0 _0421_
rlabel metal1 5888 7990 5888 7990 0 _0422_
rlabel metal2 5842 8330 5842 8330 0 _0423_
rlabel metal1 5382 6120 5382 6120 0 _0424_
rlabel metal1 5060 5882 5060 5882 0 _0425_
rlabel metal2 7498 5780 7498 5780 0 _0426_
rlabel metal2 5750 5542 5750 5542 0 _0427_
rlabel metal1 8280 5814 8280 5814 0 _0428_
rlabel metal1 8234 5338 8234 5338 0 _0429_
rlabel metal1 8326 6290 8326 6290 0 _0430_
rlabel metal1 9552 6358 9552 6358 0 _0431_
rlabel metal1 8970 9044 8970 9044 0 _0432_
rlabel metal1 12834 19176 12834 19176 0 _0433_
rlabel via2 13478 20451 13478 20451 0 _0434_
rlabel metal2 12834 21556 12834 21556 0 _0435_
rlabel metal2 13202 21148 13202 21148 0 _0436_
rlabel metal1 11362 22542 11362 22542 0 _0437_
rlabel metal2 11730 21726 11730 21726 0 _0438_
rlabel metal1 3450 14416 3450 14416 0 _0439_
rlabel metal1 2990 15130 2990 15130 0 _0440_
rlabel metal1 2162 15402 2162 15402 0 _0441_
rlabel metal1 2553 15470 2553 15470 0 _0442_
rlabel metal1 2422 15402 2422 15402 0 _0443_
rlabel metal2 1426 11934 1426 11934 0 _0444_
rlabel metal1 3358 13940 3358 13940 0 _0445_
rlabel metal2 3358 13430 3358 13430 0 _0446_
rlabel metal1 2024 11866 2024 11866 0 _0447_
rlabel metal1 2576 12206 2576 12206 0 _0448_
rlabel metal1 3036 11866 3036 11866 0 _0449_
rlabel metal1 3864 12818 3864 12818 0 _0450_
rlabel via1 3439 12138 3439 12138 0 _0451_
rlabel metal1 7971 10982 7971 10982 0 _0452_
rlabel metal2 4278 11169 4278 11169 0 _0453_
rlabel metal1 4058 11050 4058 11050 0 _0454_
rlabel metal1 5596 10710 5596 10710 0 _0455_
rlabel metal2 8326 11662 8326 11662 0 _0456_
rlabel metal1 7636 11118 7636 11118 0 _0457_
rlabel via1 7414 11050 7414 11050 0 _0458_
rlabel metal1 9246 13294 9246 13294 0 _0459_
rlabel metal1 8602 12172 8602 12172 0 _0460_
rlabel metal1 8664 11050 8664 11050 0 _0461_
rlabel via1 8978 12886 8978 12886 0 _0462_
rlabel metal2 10074 13702 10074 13702 0 _0463_
rlabel metal1 9890 13872 9890 13872 0 _0464_
rlabel metal1 9844 13974 9844 13974 0 _0465_
rlabel metal1 22310 17306 22310 17306 0 _0466_
rlabel metal1 24656 17714 24656 17714 0 _0467_
rlabel metal1 24334 15946 24334 15946 0 _0468_
rlabel metal2 13110 12070 13110 12070 0 _0469_
rlabel metal2 19366 20196 19366 20196 0 _0470_
rlabel metal1 18354 20502 18354 20502 0 _0471_
rlabel metal1 18676 20502 18676 20502 0 _0472_
rlabel metal1 20930 21930 20930 21930 0 _0473_
rlabel metal1 20838 20570 20838 20570 0 _0474_
rlabel metal2 21022 21165 21022 21165 0 _0475_
rlabel metal1 20562 19822 20562 19822 0 _0476_
rlabel metal2 19090 19686 19090 19686 0 _0477_
rlabel metal1 19688 22406 19688 22406 0 _0478_
rlabel metal2 21850 18428 21850 18428 0 _0479_
rlabel metal1 18814 18258 18814 18258 0 _0480_
rlabel metal1 20102 17238 20102 17238 0 _0481_
rlabel metal1 21068 17170 21068 17170 0 _0482_
rlabel metal1 21528 18258 21528 18258 0 _0483_
rlabel metal2 20516 18258 20516 18258 0 _0484_
rlabel metal1 20240 16558 20240 16558 0 _0485_
rlabel metal2 21114 16762 21114 16762 0 _0486_
rlabel metal1 20608 16626 20608 16626 0 _0487_
rlabel metal2 21942 17000 21942 17000 0 _0488_
rlabel metal1 19458 17102 19458 17102 0 _0489_
rlabel metal1 21942 21862 21942 21862 0 _0490_
rlabel metal1 17204 20910 17204 20910 0 _0491_
rlabel metal1 20930 23120 20930 23120 0 _0492_
rlabel metal1 22954 21658 22954 21658 0 _0493_
rlabel metal1 22678 20910 22678 20910 0 _0494_
rlabel metal1 23690 21114 23690 21114 0 _0495_
rlabel metal1 22586 20978 22586 20978 0 _0496_
rlabel metal1 22724 19958 22724 19958 0 _0497_
rlabel metal1 23782 20570 23782 20570 0 _0498_
rlabel metal1 22034 19312 22034 19312 0 _0499_
rlabel metal2 22494 19686 22494 19686 0 _0500_
rlabel metal1 23276 18394 23276 18394 0 _0501_
rlabel metal1 24104 18938 24104 18938 0 _0502_
rlabel metal2 21666 18428 21666 18428 0 _0503_
rlabel metal1 23598 16660 23598 16660 0 _0504_
rlabel metal2 22126 15572 22126 15572 0 _0505_
rlabel metal1 23322 16218 23322 16218 0 _0506_
rlabel via2 20378 20893 20378 20893 0 _0507_
rlabel metal2 20746 20978 20746 20978 0 _0508_
rlabel metal2 20194 21114 20194 21114 0 _0509_
rlabel metal2 20470 15793 20470 15793 0 _0510_
rlabel metal2 21942 15521 21942 15521 0 _0511_
rlabel metal2 23782 15368 23782 15368 0 _0512_
rlabel metal2 19458 23562 19458 23562 0 _0513_
rlabel metal1 13662 8296 13662 8296 0 _0514_
rlabel metal1 12972 11118 12972 11118 0 _0515_
rlabel metal1 12236 11050 12236 11050 0 _0516_
rlabel metal1 17250 21012 17250 21012 0 _0517_
rlabel metal2 14674 9690 14674 9690 0 _0518_
rlabel metal1 14812 11322 14812 11322 0 _0519_
rlabel metal1 17296 24106 17296 24106 0 _0520_
rlabel metal1 18262 22474 18262 22474 0 _0521_
rlabel metal1 14030 11628 14030 11628 0 _0522_
rlabel metal1 17434 21998 17434 21998 0 _0523_
rlabel metal2 23598 18326 23598 18326 0 _0524_
rlabel metal1 22954 16048 22954 16048 0 _0525_
rlabel metal1 24058 15878 24058 15878 0 _0526_
rlabel metal3 751 18428 751 18428 0 b0
rlabel metal3 751 21148 751 21148 0 b1
rlabel metal1 13294 14008 13294 14008 0 clk
rlabel metal1 16928 17646 16928 17646 0 clknet_0_clk
rlabel metal1 2070 4658 2070 4658 0 clknet_4_0_0_clk
rlabel metal2 19090 5984 19090 5984 0 clknet_4_10_0_clk
rlabel metal1 21022 9010 21022 9010 0 clknet_4_11_0_clk
rlabel metal1 17250 17238 17250 17238 0 clknet_4_12_0_clk
rlabel metal1 15318 21522 15318 21522 0 clknet_4_13_0_clk
rlabel metal1 24242 13294 24242 13294 0 clknet_4_14_0_clk
rlabel metal1 23690 21522 23690 21522 0 clknet_4_15_0_clk
rlabel metal1 1702 11764 1702 11764 0 clknet_4_1_0_clk
rlabel metal2 8786 6256 8786 6256 0 clknet_4_2_0_clk
rlabel metal1 11178 12750 11178 12750 0 clknet_4_3_0_clk
rlabel metal1 1978 17646 1978 17646 0 clknet_4_4_0_clk
rlabel metal1 7682 21556 7682 21556 0 clknet_4_5_0_clk
rlabel metal1 13662 15028 13662 15028 0 clknet_4_6_0_clk
rlabel metal2 12926 20094 12926 20094 0 clknet_4_7_0_clk
rlabel metal2 18170 4624 18170 4624 0 clknet_4_8_0_clk
rlabel metal2 14766 11968 14766 11968 0 clknet_4_9_0_clk
rlabel metal2 25898 22797 25898 22797 0 compr
rlabel metal1 12742 14416 12742 14416 0 control.baud_clk
rlabel metal1 2346 14824 2346 14824 0 control.baud_rate_gen.count\[0\]
rlabel metal1 9292 12614 9292 12614 0 control.baud_rate_gen.count\[10\]
rlabel metal1 8970 13226 8970 13226 0 control.baud_rate_gen.count\[11\]
rlabel metal1 8510 14926 8510 14926 0 control.baud_rate_gen.count\[12\]
rlabel metal1 3772 15402 3772 15402 0 control.baud_rate_gen.count\[1\]
rlabel metal1 3910 15878 3910 15878 0 control.baud_rate_gen.count\[2\]
rlabel metal1 4784 14586 4784 14586 0 control.baud_rate_gen.count\[3\]
rlabel metal1 4600 11866 4600 11866 0 control.baud_rate_gen.count\[4\]
rlabel metal2 4738 12172 4738 12172 0 control.baud_rate_gen.count\[5\]
rlabel metal2 3634 11186 3634 11186 0 control.baud_rate_gen.count\[6\]
rlabel metal1 5704 12886 5704 12886 0 control.baud_rate_gen.count\[7\]
rlabel metal1 7958 11662 7958 11662 0 control.baud_rate_gen.count\[8\]
rlabel metal1 8418 11866 8418 11866 0 control.baud_rate_gen.count\[9\]
rlabel via1 10253 14994 10253 14994 0 control.baud_rate_gen.n805_o
rlabel metal1 16836 21998 16836 21998 0 control.n576_q\[0\]
rlabel metal1 16560 21930 16560 21930 0 control.n576_q\[1\]
rlabel metal1 16836 22066 16836 22066 0 control.n576_q\[2\]
rlabel metal1 15042 22950 15042 22950 0 control.n579_q
rlabel metal1 21942 23052 21942 23052 0 control.n588_o
rlabel metal1 25116 22610 25116 22610 0 control.n598_o
rlabel metal1 24334 21658 24334 21658 0 control.n600_o
rlabel metal1 25300 19482 25300 19482 0 control.n602_o
rlabel metal2 25530 16252 25530 16252 0 control.n604_o
rlabel metal1 25484 18734 25484 18734 0 control.n606_o
rlabel metal2 25162 17476 25162 17476 0 control.n608_o
rlabel metal1 25760 20434 25760 20434 0 control.n610_o
rlabel metal1 24978 15572 24978 15572 0 control.n612_o
rlabel metal1 17066 20570 17066 20570 0 control.n633_o
rlabel metal2 19274 19754 19274 19754 0 control.n635_o
rlabel metal2 18354 16660 18354 16660 0 control.n637_o
rlabel metal2 16882 17340 16882 17340 0 control.n639_o
rlabel metal2 18722 15674 18722 15674 0 control.n641_o
rlabel metal2 20286 15640 20286 15640 0 control.n643_o
rlabel metal1 18446 16762 18446 16762 0 control.n645_o
rlabel metal1 17296 20026 17296 20026 0 control.n647_o
rlabel metal1 21160 22134 21160 22134 0 control.n651_o
rlabel metal2 20194 23562 20194 23562 0 control.n653_o
rlabel metal3 26182 21828 26182 21828 0 dac[0]
rlabel metal2 25438 21505 25438 21505 0 dac[1]
rlabel metal2 24150 19737 24150 19737 0 dac[2]
rlabel via2 25806 17051 25806 17051 0 dac[3]
rlabel metal2 25438 18751 25438 18751 0 dac[4]
rlabel metal2 25806 17901 25806 17901 0 dac[5]
rlabel metal1 25898 21862 25898 21862 0 dac[6]
rlabel metal2 25438 15181 25438 15181 0 dac[7]
rlabel metal2 11638 1520 11638 1520 0 dac_coupl
rlabel metal3 751 15708 751 15708 0 m0
rlabel metal3 1096 15028 1096 15028 0 m1
rlabel metal2 18998 10438 18998 10438 0 n119_q\[0\]
rlabel metal1 19964 9486 19964 9486 0 n119_q\[1\]
rlabel metal1 18814 12138 18814 12138 0 n119_q\[2\]
rlabel metal1 14858 22746 14858 22746 0 n120_q
rlabel metal2 15410 17986 15410 17986 0 n126_q\[0\]
rlabel metal1 18400 13498 18400 13498 0 n126_q\[1\]
rlabel metal1 18354 17238 18354 17238 0 n126_q\[2\]
rlabel metal1 16192 14042 16192 14042 0 n126_q\[3\]
rlabel metal1 18722 14586 18722 14586 0 n126_q\[4\]
rlabel metal1 14536 14790 14536 14790 0 n126_q\[5\]
rlabel metal2 18538 14722 18538 14722 0 n126_q\[6\]
rlabel metal2 17158 16558 17158 16558 0 n126_q\[7\]
rlabel metal2 13294 17204 13294 17204 0 n127_q
rlabel metal2 6854 17799 6854 17799 0 net1
rlabel metal1 23874 19482 23874 19482 0 net10
rlabel metal2 13754 8874 13754 8874 0 net100
rlabel metal2 12282 10438 12282 10438 0 net101
rlabel metal1 15456 13158 15456 13158 0 net102
rlabel metal2 16054 17884 16054 17884 0 net103
rlabel metal1 17296 14994 17296 14994 0 net104
rlabel metal2 13570 13770 13570 13770 0 net105
rlabel metal2 12926 15980 12926 15980 0 net106
rlabel metal1 18768 12954 18768 12954 0 net107
rlabel metal2 19826 14144 19826 14144 0 net108
rlabel metal2 12466 7582 12466 7582 0 net109
rlabel metal2 24794 16524 24794 16524 0 net11
rlabel metal1 19320 17170 19320 17170 0 net110
rlabel metal1 15732 17714 15732 17714 0 net111
rlabel metal1 17342 20774 17342 20774 0 net112
rlabel metal1 20102 16762 20102 16762 0 net113
rlabel metal1 15778 15130 15778 15130 0 net114
rlabel metal2 19274 11526 19274 11526 0 net115
rlabel metal1 13662 16082 13662 16082 0 net116
rlabel metal1 21942 16592 21942 16592 0 net117
rlabel metal2 10994 23868 10994 23868 0 net118
rlabel metal2 12190 23494 12190 23494 0 net119
rlabel metal1 25300 18258 25300 18258 0 net12
rlabel metal1 9660 6766 9660 6766 0 net120
rlabel metal1 8924 6426 8924 6426 0 net121
rlabel metal2 16054 22780 16054 22780 0 net122
rlabel metal1 15512 23086 15512 23086 0 net123
rlabel metal2 11914 21760 11914 21760 0 net124
rlabel metal1 17894 22066 17894 22066 0 net125
rlabel metal1 14628 21862 14628 21862 0 net126
rlabel metal1 10488 9350 10488 9350 0 net127
rlabel metal2 12558 8364 12558 8364 0 net128
rlabel metal2 12374 8296 12374 8296 0 net129
rlabel metal1 25530 17306 25530 17306 0 net13
rlabel metal1 17940 12138 17940 12138 0 net130
rlabel metal2 13294 24480 13294 24480 0 net131
rlabel metal1 13616 20570 13616 20570 0 net132
rlabel metal1 20056 15470 20056 15470 0 net133
rlabel metal1 21160 19822 21160 19822 0 net134
rlabel metal1 12466 23120 12466 23120 0 net135
rlabel metal2 18722 23052 18722 23052 0 net136
rlabel metal1 13754 19788 13754 19788 0 net137
rlabel metal1 19872 9962 19872 9962 0 net138
rlabel metal1 25300 20570 25300 20570 0 net14
rlabel metal1 25208 15130 25208 15130 0 net15
rlabel metal1 11960 5542 11960 5542 0 net16
rlabel metal1 20700 6630 20700 6630 0 net17
rlabel metal2 23966 12988 23966 12988 0 net18
rlabel metal2 25254 6188 25254 6188 0 net19
rlabel metal2 3266 21148 3266 21148 0 net2
rlabel metal2 20562 6596 20562 6596 0 net20
rlabel metal1 25760 14246 25760 14246 0 net21
rlabel metal1 21390 2482 21390 2482 0 net22
rlabel metal1 22862 4046 22862 4046 0 net23
rlabel metal1 22862 6664 22862 6664 0 net24
rlabel metal1 16008 2414 16008 2414 0 net25
rlabel metal1 18216 3094 18216 3094 0 net26
rlabel metal1 19964 3978 19964 3978 0 net27
rlabel metal1 15457 3026 15457 3026 0 net28
rlabel metal2 18630 2516 18630 2516 0 net29
rlabel metal1 20470 21590 20470 21590 0 net3
rlabel metal2 17250 4012 17250 4012 0 net30
rlabel metal2 17802 2587 17802 2587 0 net31
rlabel metal1 20516 5202 20516 5202 0 net32
rlabel metal1 25116 5610 25116 5610 0 net33
rlabel metal1 23322 3910 23322 3910 0 net34
rlabel metal2 23874 3519 23874 3519 0 net35
rlabel metal1 25438 5338 25438 5338 0 net36
rlabel metal1 23000 2414 23000 2414 0 net37
rlabel metal1 24564 6086 24564 6086 0 net38
rlabel metal1 21298 2346 21298 2346 0 net39
rlabel metal2 1610 16320 1610 16320 0 net4
rlabel metal1 20884 4590 20884 4590 0 net40
rlabel metal1 25070 8330 25070 8330 0 net41
rlabel metal1 25070 11594 25070 11594 0 net42
rlabel metal1 25208 10438 25208 10438 0 net43
rlabel metal1 25208 7514 25208 7514 0 net44
rlabel metal1 25438 12104 25438 12104 0 net45
rlabel metal1 25668 7378 25668 7378 0 net46
rlabel metal1 24288 11526 24288 11526 0 net47
rlabel metal1 23138 8942 23138 8942 0 net48
rlabel metal1 13708 2414 13708 2414 0 net49
rlabel metal1 1702 15674 1702 15674 0 net5
rlabel metal1 21298 12104 21298 12104 0 net50
rlabel metal2 21390 12257 21390 12257 0 net51
rlabel metal1 14306 2414 14306 2414 0 net52
rlabel metal1 21666 14450 21666 14450 0 net53
rlabel via1 14306 6086 14306 6086 0 net54
rlabel metal1 21712 13770 21712 13770 0 net55
rlabel metal1 16698 2414 16698 2414 0 net56
rlabel metal2 13202 25806 13202 25806 0 net57
rlabel metal2 2530 5984 2530 5984 0 net58
rlabel metal1 2484 20434 2484 20434 0 net59
rlabel metal1 12466 13940 12466 13940 0 net6
rlabel metal2 2530 12121 2530 12121 0 net60
rlabel metal1 8700 13872 8700 13872 0 net61
rlabel metal1 2530 21998 2530 21998 0 net62
rlabel via1 13390 14994 13390 14994 0 net63
rlabel metal1 20654 20332 20654 20332 0 net64
rlabel metal1 16146 17748 16146 17748 0 net65
rlabel metal1 23644 12886 23644 12886 0 net66
rlabel metal1 19090 20400 19090 20400 0 net67
rlabel metal2 2714 21216 2714 21216 0 net68
rlabel metal1 7866 18190 7866 18190 0 net69
rlabel metal1 10534 2618 10534 2618 0 net7
rlabel metal2 15134 5440 15134 5440 0 net70
rlabel metal1 6670 18768 6670 18768 0 net71
rlabel via1 6670 7854 6670 7854 0 net72
rlabel metal1 13938 5134 13938 5134 0 net73
rlabel metal1 21850 4794 21850 4794 0 net74
rlabel metal2 21482 7055 21482 7055 0 net75
rlabel metal1 20746 14348 20746 14348 0 net76
rlabel metal1 21206 13294 21206 13294 0 net77
rlabel metal2 19274 18496 19274 18496 0 net78
rlabel metal1 6256 20910 6256 20910 0 net79
rlabel metal2 25622 22780 25622 22780 0 net8
rlabel metal1 4094 7310 4094 7310 0 net80
rlabel metal1 6716 8942 6716 8942 0 net81
rlabel metal1 13887 22678 13887 22678 0 net82
rlabel metal1 9844 7718 9844 7718 0 net83
rlabel metal2 18630 18428 18630 18428 0 net84
rlabel metal2 18998 14144 18998 14144 0 net85
rlabel metal1 25024 19754 25024 19754 0 net86
rlabel metal1 25024 17578 25024 17578 0 net87
rlabel metal1 25024 18666 25024 18666 0 net88
rlabel metal1 24840 22542 24840 22542 0 net89
rlabel metal2 23690 21658 23690 21658 0 net9
rlabel metal1 24702 20502 24702 20502 0 net90
rlabel metal1 15134 18598 15134 18598 0 net91
rlabel metal1 11523 6290 11523 6290 0 net92
rlabel metal1 24012 15130 24012 15130 0 net93
rlabel metal1 24564 20910 24564 20910 0 net94
rlabel metal2 15318 19788 15318 19788 0 net95
rlabel metal1 24380 16218 24380 16218 0 net96
rlabel metal2 18722 20604 18722 20604 0 net97
rlabel metal1 10764 22066 10764 22066 0 net98
rlabel metal1 12742 17000 12742 17000 0 net99
rlabel metal2 20654 1520 20654 1520 0 reg0[0]
rlabel via2 25806 12971 25806 12971 0 reg0[1]
rlabel via2 25806 2805 25806 2805 0 reg0[2]
rlabel metal2 25806 3417 25806 3417 0 reg0[3]
rlabel metal2 25806 15793 25806 15793 0 reg0[4]
rlabel metal2 21298 1690 21298 1690 0 reg0[5]
rlabel metal2 25438 4063 25438 4063 0 reg0[6]
rlabel metal2 25438 6749 25438 6749 0 reg0[7]
rlabel metal2 15502 1520 15502 1520 0 reg1[0]
rlabel metal2 18078 1520 18078 1520 0 reg1[1]
rlabel metal2 19366 959 19366 959 0 reg1[2]
rlabel metal2 14858 1520 14858 1520 0 reg1[3]
rlabel metal2 18722 1656 18722 1656 0 reg1[4]
rlabel metal2 16790 1520 16790 1520 0 reg1[5]
rlabel metal2 17434 1520 17434 1520 0 reg1[6]
rlabel metal2 20010 1520 20010 1520 0 reg1[7]
rlabel metal2 25806 4403 25806 4403 0 reg2[0]
rlabel metal2 24518 1520 24518 1520 0 reg2[1]
rlabel metal2 23874 1520 23874 1520 0 reg2[2]
rlabel metal2 25806 5423 25806 5423 0 reg2[3]
rlabel metal2 22586 1520 22586 1520 0 reg2[4]
rlabel metal2 25806 6035 25806 6035 0 reg2[5]
rlabel metal2 21942 1588 21942 1588 0 reg2[6]
rlabel metal2 23230 1520 23230 1520 0 reg2[7]
rlabel metal2 25806 8857 25806 8857 0 reg3[0]
rlabel via2 25806 10251 25806 10251 0 reg3[1]
rlabel metal2 25806 10863 25806 10863 0 reg3[2]
rlabel metal2 25806 7089 25806 7089 0 reg3[3]
rlabel metal2 25806 12087 25806 12087 0 reg3[4]
rlabel metal1 25990 7514 25990 7514 0 reg3[5]
rlabel metal2 25806 11475 25806 11475 0 reg3[6]
rlabel metal2 25438 9741 25438 9741 0 reg3[7]
rlabel metal2 12926 1520 12926 1520 0 reg4[0]
rlabel metal2 25806 14195 25806 14195 0 reg4[1]
rlabel metal2 25438 13855 25438 13855 0 reg4[2]
rlabel metal2 14214 1520 14214 1520 0 reg4[3]
rlabel metal1 25944 15674 25944 15674 0 reg4[4]
rlabel metal2 13570 1520 13570 1520 0 reg4[5]
rlabel metal2 25806 18955 25806 18955 0 reg4[6]
rlabel metal2 16146 1520 16146 1520 0 reg4[7]
rlabel metal2 12282 1588 12282 1588 0 rst
rlabel metal2 10350 1588 10350 1588 0 rx
rlabel metal1 13018 27098 13018 27098 0 tx
rlabel metal2 9614 8908 9614 8908 0 uart_receive.baud_clk
rlabel metal1 11040 8398 11040 8398 0 uart_receive.baud_clk2
rlabel metal1 13754 9010 13754 9010 0 uart_receive.baud_clk3
rlabel metal2 2714 5440 2714 5440 0 uart_receive.baud_rate_gen.count\[0\]
rlabel metal1 8602 7378 8602 7378 0 uart_receive.baud_rate_gen.count\[10\]
rlabel metal2 7866 7174 7866 7174 0 uart_receive.baud_rate_gen.count\[11\]
rlabel metal2 2622 5848 2622 5848 0 uart_receive.baud_rate_gen.count\[1\]
rlabel metal2 2162 6494 2162 6494 0 uart_receive.baud_rate_gen.count\[2\]
rlabel metal1 3358 7174 3358 7174 0 uart_receive.baud_rate_gen.count\[3\]
rlabel metal1 5382 8976 5382 8976 0 uart_receive.baud_rate_gen.count\[4\]
rlabel metal2 5474 9044 5474 9044 0 uart_receive.baud_rate_gen.count\[5\]
rlabel via2 5658 8891 5658 8891 0 uart_receive.baud_rate_gen.count\[6\]
rlabel metal2 6900 7854 6900 7854 0 uart_receive.baud_rate_gen.count\[7\]
rlabel metal1 6624 5814 6624 5814 0 uart_receive.baud_rate_gen.count\[8\]
rlabel metal1 8694 7174 8694 7174 0 uart_receive.baud_rate_gen.count\[9\]
rlabel metal1 11178 7514 11178 7514 0 uart_receive.n328_o\[0\]
rlabel via1 11357 6766 11357 6766 0 uart_receive.n328_o\[1\]
rlabel metal1 8234 7956 8234 7956 0 uart_receive.n345_q
rlabel metal1 12834 8262 12834 8262 0 uart_receive.n346_q\[0\]
rlabel metal1 13386 8500 13386 8500 0 uart_receive.n346_q\[1\]
rlabel metal1 12696 11866 12696 11866 0 uart_receive.n352_o
rlabel metal1 13202 12614 13202 12614 0 uart_receive.n354_o
rlabel metal2 12926 9248 12926 9248 0 uart_receive.n360_o
rlabel metal2 18446 10302 18446 10302 0 uart_receive.n370_o
rlabel metal1 21068 12818 21068 12818 0 uart_receive.n372_o
rlabel metal1 19458 3502 19458 3502 0 uart_receive.n374_o
rlabel metal2 21758 6595 21758 6595 0 uart_receive.n376_o
rlabel metal1 16422 9452 16422 9452 0 uart_receive.n378_o
rlabel metal2 19182 7327 19182 7327 0 uart_receive.n380_o
rlabel via2 16974 3043 16974 3043 0 uart_receive.n382_o
rlabel metal1 20562 8942 20562 8942 0 uart_receive.n384_o
rlabel metal2 13202 22882 13202 22882 0 uart_transmit.baud_clk
rlabel metal2 4002 17952 4002 17952 0 uart_transmit.baud_rate_gen.count\[0\]
rlabel metal1 8188 18598 8188 18598 0 uart_transmit.baud_rate_gen.count\[10\]
rlabel metal2 8970 18258 8970 18258 0 uart_transmit.baud_rate_gen.count\[11\]
rlabel metal2 6486 18496 6486 18496 0 uart_transmit.baud_rate_gen.count\[12\]
rlabel metal2 2254 18870 2254 18870 0 uart_transmit.baud_rate_gen.count\[1\]
rlabel metal1 3220 20502 3220 20502 0 uart_transmit.baud_rate_gen.count\[2\]
rlabel metal1 3496 20910 3496 20910 0 uart_transmit.baud_rate_gen.count\[3\]
rlabel metal1 5336 21930 5336 21930 0 uart_transmit.baud_rate_gen.count\[4\]
rlabel metal1 5428 21862 5428 21862 0 uart_transmit.baud_rate_gen.count\[5\]
rlabel metal1 5750 20978 5750 20978 0 uart_transmit.baud_rate_gen.count\[6\]
rlabel metal1 6854 20978 6854 20978 0 uart_transmit.baud_rate_gen.count\[7\]
rlabel metal1 7498 18224 7498 18224 0 uart_transmit.baud_rate_gen.count\[8\]
rlabel metal2 7406 19754 7406 19754 0 uart_transmit.baud_rate_gen.count\[9\]
rlabel metal2 13570 21828 13570 21828 0 uart_transmit.n167_o
rlabel metal2 9430 24310 9430 24310 0 uart_transmit.n224_q
rlabel metal2 12466 23256 12466 23256 0 uart_transmit.n226_q\[0\]
rlabel metal2 13386 23018 13386 23018 0 uart_transmit.n226_q\[1\]
rlabel metal2 14398 20740 14398 20740 0 uart_transmit.n227_q\[0\]
rlabel metal1 14214 20468 14214 20468 0 uart_transmit.n227_q\[1\]
rlabel metal1 14122 19278 14122 19278 0 uart_transmit.n227_q\[2\]
rlabel metal1 11362 21998 11362 21998 0 uart_transmit.n227_q\[3\]
rlabel metal2 12558 21284 12558 21284 0 uart_transmit.n227_q\[4\]
rlabel metal1 14352 20026 14352 20026 0 uart_transmit.n231_o
rlabel metal2 12926 17544 12926 17544 0 uart_transmit.n232_o
rlabel metal1 12696 16218 12696 16218 0 uart_transmit.n233_o
rlabel metal1 14398 16116 14398 16116 0 uart_transmit.n234_o
rlabel metal2 14122 18598 14122 18598 0 uart_transmit.n235_o
rlabel metal1 14352 16966 14352 16966 0 uart_transmit.n236_o
rlabel metal2 14490 18564 14490 18564 0 uart_transmit.n237_o
<< properties >>
string FIXED_BBOX 0 0 27332 29476
<< end >>
