magic
tech sky130A
magscale 1 2
timestamp 1730928274
<< locali >>
rect -60 1340 1080 1440
rect 260 1280 760 1340
rect 2300 0 2800 40
rect 1160 -100 4100 0
<< metal1 >>
rect -60 1140 740 1240
rect 1020 1160 3960 1260
rect -60 180 40 1140
rect 140 980 200 1000
rect 140 880 200 920
rect 140 800 200 820
rect 330 980 390 1000
rect 330 880 390 920
rect 330 800 390 820
rect 520 980 580 1000
rect 520 880 580 920
rect 520 800 580 820
rect 710 980 770 1000
rect 710 880 770 920
rect 710 800 770 820
rect 230 480 290 500
rect 230 380 290 420
rect 230 300 290 320
rect 420 480 480 500
rect 420 380 480 420
rect 420 300 480 320
rect 620 480 680 500
rect 620 380 680 420
rect 620 300 680 320
rect 810 480 870 500
rect 810 380 870 420
rect 810 300 870 320
rect 1020 180 1120 1160
rect 1240 980 1300 1000
rect 1240 880 1300 920
rect 1240 800 1300 820
rect 1490 980 1550 1000
rect 1490 880 1550 920
rect 1490 800 1550 820
rect 1750 980 1810 1000
rect 1750 880 1810 920
rect 1750 800 1810 820
rect 2000 980 2060 1000
rect 2000 880 2060 920
rect 2000 800 2060 820
rect 2260 980 2320 1000
rect 2260 880 2320 920
rect 2260 800 2320 820
rect 2520 980 2580 1000
rect 2520 880 2580 920
rect 2520 800 2580 820
rect 2770 980 2830 1000
rect 2770 880 2830 920
rect 2770 800 2830 820
rect 3030 980 3090 1000
rect 3030 880 3090 920
rect 3030 800 3090 820
rect 3280 980 3340 1000
rect 3280 880 3340 920
rect 3280 800 3340 820
rect 3540 980 3600 1000
rect 3540 880 3600 920
rect 3540 800 3600 820
rect 3800 980 3860 1000
rect 3800 880 3860 920
rect 3800 800 3860 820
rect 1360 480 1420 500
rect 1360 380 1420 420
rect 1360 300 1420 320
rect 1620 480 1680 500
rect 1620 380 1680 420
rect 1620 300 1680 320
rect 1880 480 1940 500
rect 1880 380 1940 420
rect 1880 300 1940 320
rect 2130 480 2190 500
rect 2130 380 2190 420
rect 2130 300 2190 320
rect 2390 480 2450 500
rect 2390 380 2450 420
rect 2390 300 2450 320
rect 2640 480 2700 500
rect 2640 380 2700 420
rect 2640 300 2700 320
rect 2900 480 2960 500
rect 2900 380 2960 420
rect 2900 300 2960 320
rect 3160 480 3220 500
rect 3160 380 3220 420
rect 3160 300 3220 320
rect 3410 480 3470 500
rect 3410 380 3470 420
rect 3410 300 3470 320
rect 3670 480 3730 500
rect 3670 380 3730 420
rect 3670 300 3730 320
rect 3930 480 3990 500
rect 3930 380 3990 420
rect 3930 300 3990 320
rect -60 80 840 180
rect 1020 80 3960 180
<< via1 >>
rect 140 920 200 980
rect 140 820 200 880
rect 330 920 390 980
rect 330 820 390 880
rect 520 920 580 980
rect 520 820 580 880
rect 710 920 770 980
rect 710 820 770 880
rect 230 420 290 480
rect 230 320 290 380
rect 420 420 480 480
rect 420 320 480 380
rect 620 420 680 480
rect 620 320 680 380
rect 810 420 870 480
rect 810 320 870 380
rect 1240 920 1300 980
rect 1240 820 1300 880
rect 1490 920 1550 980
rect 1490 820 1550 880
rect 1750 920 1810 980
rect 1750 820 1810 880
rect 2000 920 2060 980
rect 2000 820 2060 880
rect 2260 920 2320 980
rect 2260 820 2320 880
rect 2520 920 2580 980
rect 2520 820 2580 880
rect 2770 920 2830 980
rect 2770 820 2830 880
rect 3030 920 3090 980
rect 3030 820 3090 880
rect 3280 920 3340 980
rect 3280 820 3340 880
rect 3540 920 3600 980
rect 3540 820 3600 880
rect 3800 920 3860 980
rect 3800 820 3860 880
rect 1360 420 1420 480
rect 1360 320 1420 380
rect 1620 420 1680 480
rect 1620 320 1680 380
rect 1880 420 1940 480
rect 1880 320 1940 380
rect 2130 420 2190 480
rect 2130 320 2190 380
rect 2390 420 2450 480
rect 2390 320 2450 380
rect 2640 420 2700 480
rect 2640 320 2700 380
rect 2900 420 2960 480
rect 2900 320 2960 380
rect 3160 420 3220 480
rect 3160 320 3220 380
rect 3410 420 3470 480
rect 3410 320 3470 380
rect 3670 420 3730 480
rect 3670 320 3730 380
rect 3930 420 3990 480
rect 3930 320 3990 380
<< metal2 >>
rect 100 980 4400 1000
rect 100 920 140 980
rect 200 920 330 980
rect 390 920 520 980
rect 580 920 710 980
rect 770 920 1240 980
rect 1300 920 1490 980
rect 1550 920 1750 980
rect 1810 920 2000 980
rect 2060 920 2260 980
rect 2320 920 2520 980
rect 2580 920 2770 980
rect 2830 920 3030 980
rect 3090 920 3280 980
rect 3340 920 3540 980
rect 3600 920 3800 980
rect 3860 920 4400 980
rect 100 880 4400 920
rect 100 820 140 880
rect 200 820 330 880
rect 390 820 520 880
rect 580 820 710 880
rect 770 820 1240 880
rect 1300 820 1490 880
rect 1550 820 1750 880
rect 1810 820 2000 880
rect 2060 820 2260 880
rect 2320 820 2520 880
rect 2580 820 2770 880
rect 2830 820 3030 880
rect 3090 820 3280 880
rect 3340 820 3540 880
rect 3600 820 3800 880
rect 3860 820 4400 880
rect 100 800 4400 820
rect 100 480 4400 500
rect 100 420 230 480
rect 290 420 420 480
rect 480 420 620 480
rect 680 420 810 480
rect 870 420 1360 480
rect 1420 420 1620 480
rect 1680 420 1880 480
rect 1940 420 2130 480
rect 2190 420 2390 480
rect 2450 420 2640 480
rect 2700 420 2900 480
rect 2960 420 3160 480
rect 3220 420 3410 480
rect 3470 420 3670 480
rect 3730 420 3930 480
rect 3990 420 4400 480
rect 100 380 4400 420
rect 100 320 230 380
rect 290 320 420 380
rect 480 320 620 380
rect 680 320 810 380
rect 870 320 1360 380
rect 1420 320 1620 380
rect 1680 320 1880 380
rect 1940 320 2130 380
rect 2190 320 2390 380
rect 2450 320 2640 380
rect 2700 320 2900 380
rect 2960 320 3160 380
rect 3220 320 3410 380
rect 3470 320 3670 380
rect 3730 320 3930 380
rect 3990 320 4400 380
rect 100 300 4400 320
use sky130_fd_pr__nfet_01v8_lvt_8AG63Z  sky130_fd_pr__nfet_01v8_lvt_8AG63Z_0
timestamp 1730928108
transform 1 0 503 0 1 660
box -503 -660 503 660
use sky130_fd_pr__pfet_01v8_lvt_MUCXQQ  sky130_fd_pr__pfet_01v8_lvt_MUCXQQ_0
timestamp 1730928108
transform 1 0 2611 0 1 669
box -1511 -669 1511 669
<< labels >>
rlabel locali 1160 -100 1260 0 1 VPWR
port 1 n
rlabel locali -60 1340 40 1440 1 VGND
port 2 n
rlabel metal1 -60 620 40 720 1 CTRL_P
port 3 n
rlabel metal1 1020 620 1120 720 1 CTRL_N
port 4 n
rlabel metal2 4200 800 4400 1000 1 X
port 5 n
rlabel metal2 4200 300 4400 500 1 Y
port 6 n
<< end >>
