* NGSPICE file created from variable_delay_parax.ext - technology: sky130A

.subckt variable_delay_parax in en_1 en_6 out en_2 en_3 en_5 en_7 en_0 en_4 VSS VDD
X0 a_20184_772# variable_delay_unit_7.out variable_delay_unit_6.out VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1 a_16354_772# variable_delay_unit_5.tristate_inverter_1.en.t2 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X2 VSS.t5 variable_delay_unit_8.tristate_inverter_1.en.t2 a_26080_352# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X3 a_19302_352# en_6.t0 VSS.t158 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X4 VDD.t58 en_1.t0 a_5444_772# VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X5 variable_delay_unit_4.in.t1 variable_delay_unit_3.in.t2 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X6 VSS.t9 variable_delay_unit_2.tristate_inverter_1.en.t2 a_8392_352# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X7 variable_delay_unit_8.out variable_delay_unit_8.forward.t2 a_25198_772# VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X8 a_20184_352# variable_delay_unit_7.out variable_delay_unit_6.out VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X9 a_16354_352# en_5.t0 VSS.t80 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X10 VDD.t54 en_1.t1 a_5444_772# VDD.t53 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X11 variable_delay_unit_3.in.t0 variable_delay_unit_2.in.t2 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X12 VDD.t131 en_0.t0 a_2496_772# VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X13 VDD.t56 en_5.t1 a_17236_772# VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X14 variable_delay_unit_4.in.t0 variable_delay_unit_3.in.t3 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 VSS.t132 variable_delay_unit_1.tristate_inverter_1.en.t2 a_5444_352# VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X16 variable_delay_unit_8.out variable_delay_unit_8.forward.t3 a_25198_352# VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X17 VSS.t122 variable_delay_unit_1.tristate_inverter_1.en.t3 a_5444_352# VSS.t121 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X18 variable_delay_unit_3.in.t1 variable_delay_unit_2.in.t3 VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X19 VSS.t38 variable_delay_unit_0.tristate_inverter_1.en.t2 a_2496_352# VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X20 VDD.t102 variable_delay_unit_2.tristate_inverter_1.en.t3 a_7510_772# VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X21 VSS.t94 variable_delay_unit_5.tristate_inverter_1.en.t3 a_17236_352# VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X22 variable_delay_unit_1.out variable_delay_unit_2.in.t4 a_4562_772# VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X23 VDD.t21 en_4.t0 a_14288_772# VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X24 a_26080_772# VSS.t163 variable_delay_unit_8.out VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X25 variable_delay_unit_6.in.t1 variable_delay_unit_5.in.t2 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X26 VDD.t157 variable_delay_unit_1.tristate_inverter_1.en.t4 a_4562_772# VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X27 VDD.t66 en_3.t0 a_11340_772# VDD.t65 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X28 variable_delay_unit_0.tristate_inverter_1.en.t1 en_0.t1 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X29 variable_delay_unit_1.out variable_delay_unit_2.in.t5 a_4562_352# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X30 VSS.t150 en_2.t0 a_7510_352# VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X31 variable_delay_unit_7.tristate_inverter_1.en.t1 en_7.t0 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X32 a_26080_352# VSS.t54 variable_delay_unit_8.out VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X33 out.t0 variable_delay_unit_1.in.t2 a_1614_772# VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X34 VSS.t45 en_1.t2 a_4562_352# VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 a_23132_772# en_7.t1 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X36 variable_delay_unit_6.in.t0 variable_delay_unit_5.in.t3 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X37 VSS.t130 variable_delay_unit_4.tristate_inverter_1.en.t2 a_14288_352# VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X38 variable_delay_unit_0.tristate_inverter_1.en.t0 en_0.t2 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X39 VSS.t86 variable_delay_unit_3.tristate_inverter_1.en.t2 a_11340_352# VSS.t85 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X40 variable_delay_unit_7.tristate_inverter_1.en.t0 en_7.t2 VSS.t119 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X41 a_23132_772# variable_delay_unit_8.out variable_delay_unit_7.out VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X42 variable_delay_unit_5.in.t1 variable_delay_unit_4.in.t2 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X43 a_20184_772# en_6.t1 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X44 VDD.t82 variable_delay_unit_4.tristate_inverter_1.en.t3 a_13406_772# VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X45 variable_delay_unit_3.out variable_delay_unit_4.in.t3 a_10458_772# VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X46 a_23132_352# variable_delay_unit_7.tristate_inverter_1.en.t2 VSS.t101 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X47 out.t1 variable_delay_unit_1.in.t3 a_1614_352# VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X48 VDD.t137 en_2.t1 a_8392_772# VDD.t136 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X49 a_23132_352# variable_delay_unit_8.out variable_delay_unit_7.out VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X50 a_25198_772# variable_delay_unit_8.tristate_inverter_1.en.t3 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X51 a_20184_352# variable_delay_unit_6.tristate_inverter_1.en.t2 VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X52 variable_delay_unit_5.in.t0 variable_delay_unit_4.in.t4 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X53 a_22250_772# variable_delay_unit_7.tristate_inverter_1.en.t3 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X54 VSS.t20 en_4.t1 a_13406_352# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X55 variable_delay_unit_3.out variable_delay_unit_4.in.t5 a_10458_352# VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X56 a_2496_772# variable_delay_unit_1.out out.t2 VDD.t151 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X57 VDD.t116 variable_delay_unit_3.tristate_inverter_1.en.t3 a_10458_772# VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X58 a_22250_772# variable_delay_unit_7.tristate_inverter_1.en.t4 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X59 VDD.t68 en_5.t2 a_17236_772# VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X60 VSS.t50 variable_delay_unit_2.tristate_inverter_1.en.t4 a_8392_352# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X61 a_25198_352# VDD.t166 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X62 a_22250_352# en_7.t3 VSS.t152 VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X63 a_2496_352# variable_delay_unit_1.out out.t3 VSS.t156 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X64 variable_delay_unit_2.out variable_delay_unit_3.in.t4 a_7510_772# VDD.t83 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X65 a_22250_352# en_7.t4 VSS.t138 VSS.t137 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X66 VSS.t92 variable_delay_unit_5.tristate_inverter_1.en.t4 a_17236_352# VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X67 VSS.t68 en_3.t1 a_10458_352# VSS.t67 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X68 variable_delay_unit_7.in.t1 variable_delay_unit_6.in.t2 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X69 VDD.t19 en_4.t2 a_14288_772# VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X70 VDD.t135 variable_delay_unit_6.tristate_inverter_1.en.t3 a_19302_772# VDD.t134 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X71 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t3 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X72 variable_delay_unit_2.out variable_delay_unit_3.in.t5 a_7510_352# VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X73 variable_delay_unit_8.tristate_inverter_1.en.t1 VDD.t78 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X74 a_26080_772# VDD.t75 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X75 variable_delay_unit_7.in.t0 variable_delay_unit_6.in.t3 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X76 VSS.t82 variable_delay_unit_4.tristate_inverter_1.en.t4 a_14288_352# VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X77 a_1614_352# en_0.t3 VSS.t31 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X78 VSS.t52 en_6.t2 a_19302_352# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X79 variable_delay_unit_5.out variable_delay_unit_6.in.t4 a_16354_772# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X80 variable_delay_unit_8.tristate_inverter_1.en.t0 VDD.t167 VSS.t76 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X81 a_5444_772# en_1.t3 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X82 a_8392_772# variable_delay_unit_3.out variable_delay_unit_2.out VDD.t145 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X83 VDD.t52 variable_delay_unit_5.tristate_inverter_1.en.t5 a_16354_772# VDD.t51 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X84 variable_delay_unit_4.out variable_delay_unit_5.in.t4 a_13406_772# VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X85 a_26080_352# variable_delay_unit_8.tristate_inverter_1.en.t4 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X86 variable_delay_unit_1.tristate_inverter_1.en.t1 en_1.t4 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X87 variable_delay_unit_5.out variable_delay_unit_6.in.t5 a_16354_352# VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X88 a_8392_352# variable_delay_unit_3.out variable_delay_unit_2.out VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X89 a_5444_352# variable_delay_unit_1.tristate_inverter_1.en.t5 VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X90 a_25198_772# variable_delay_unit_8.tristate_inverter_1.en.t5 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X91 VSS.t13 en_5.t3 a_16354_352# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X92 variable_delay_unit_4.out variable_delay_unit_5.in.t5 a_13406_352# VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X93 a_5444_772# variable_delay_unit_2.out variable_delay_unit_1.out VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X94 variable_delay_unit_1.tristate_inverter_1.en.t0 en_1.t5 VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X95 a_2496_772# en_0.t4 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X96 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en.t5 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X97 a_25198_352# VDD.t168 VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X98 a_5444_352# variable_delay_unit_2.out variable_delay_unit_1.out VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X99 a_2496_352# variable_delay_unit_0.tristate_inverter_1.en.t4 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X100 a_7510_352# en_2.t2 VSS.t146 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X101 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t6 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X102 a_11340_772# en_3.t2 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X103 a_14288_772# variable_delay_unit_5.out variable_delay_unit_4.out VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X104 VDD.t128 en_7.t5 a_23132_772# VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X105 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t5 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X106 variable_delay_unit_3.tristate_inverter_1.en.t1 en_3.t3 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X107 a_11340_772# variable_delay_unit_4.out variable_delay_unit_3.out VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X108 a_4562_352# en_1.t6 VSS.t58 VSS.t57 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X109 VSS.t134 variable_delay_unit_7.tristate_inverter_1.en.t5 a_23132_352# VSS.t133 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X110 variable_delay_unit_6.out variable_delay_unit_7.in.t2 a_19302_772# VDD.t164 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X111 a_14288_352# variable_delay_unit_5.out variable_delay_unit_4.out VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X112 a_1614_352# en_0.t5 VSS.t107 VSS.t106 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X113 variable_delay_unit_3.tristate_inverter_1.en.t0 en_3.t4 VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X114 a_11340_352# variable_delay_unit_3.tristate_inverter_1.en.t4 VSS.t128 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X115 variable_delay_unit_1.in.t0 in.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X116 variable_delay_unit_8.in.t1 variable_delay_unit_7.in.t3 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X117 VDD.t17 en_6.t3 a_20184_772# VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X118 a_11340_352# variable_delay_unit_4.out variable_delay_unit_3.out VSS.t104 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X119 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en.t5 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X120 variable_delay_unit_2.tristate_inverter_1.en.t1 en_2.t3 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X121 variable_delay_unit_6.out variable_delay_unit_7.in.t4 a_19302_352# VSS.t154 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X122 a_8392_772# en_2.t4 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X123 variable_delay_unit_1.in.t1 in.t1 VSS.t162 VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X124 variable_delay_unit_8.in.t0 variable_delay_unit_7.in.t5 VSS.t99 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X125 VSS.t26 variable_delay_unit_6.tristate_inverter_1.en.t4 a_20184_352# VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X126 variable_delay_unit_2.tristate_inverter_1.en.t0 en_2.t5 VSS.t160 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X127 a_13406_352# en_4.t3 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X128 a_17236_772# en_5.t4 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X129 a_10458_772# variable_delay_unit_3.tristate_inverter_1.en.t5 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X130 a_8392_352# variable_delay_unit_2.tristate_inverter_1.en.t6 VSS.t60 VSS.t59 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X131 variable_delay_unit_5.tristate_inverter_1.en.t1 en_5.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X132 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en.t7 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X133 a_17236_352# variable_delay_unit_5.tristate_inverter_1.en.t6 VSS.t90 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X134 a_10458_352# en_3.t5 VSS.t142 VSS.t141 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X135 variable_delay_unit_5.tristate_inverter_1.en.t0 en_5.t6 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X136 a_17236_772# variable_delay_unit_6.out variable_delay_unit_5.out VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X137 a_14288_772# en_4.t4 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X138 a_19302_772# variable_delay_unit_6.tristate_inverter_1.en.t5 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X139 a_7510_352# en_2.t6 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X140 variable_delay_unit_4.tristate_inverter_1.en.t1 en_4.t5 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X141 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t7 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X142 VDD.t74 VDD.t72 a_26080_772# VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X143 VDD.t126 en_7.t6 a_23132_772# VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X144 a_17236_352# variable_delay_unit_6.out variable_delay_unit_5.out VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X145 a_19302_352# en_6.t4 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X146 a_14288_352# variable_delay_unit_4.tristate_inverter_1.en.t6 VSS.t111 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X147 variable_delay_unit_4.tristate_inverter_1.en.t0 en_4.t6 VSS.t126 VSS.t125 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X148 a_16354_772# variable_delay_unit_5.tristate_inverter_1.en.t7 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X149 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en.t7 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X150 VSS.t1 variable_delay_unit_8.tristate_inverter_1.en.t6 a_26080_352# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X151 a_4562_352# en_1.t7 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X152 VSS.t109 variable_delay_unit_7.tristate_inverter_1.en.t6 a_23132_352# VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X153 variable_delay_unit_8.forward.t1 variable_delay_unit_8.in.t2 VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X154 VDD.t15 variable_delay_unit_8.tristate_inverter_1.en.t7 a_25198_772# VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X155 a_16354_352# en_5.t7 VSS.t41 VSS.t40 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X156 VDD.t91 en_6.t5 a_20184_772# VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X157 variable_delay_unit_7.out variable_delay_unit_8.in.t3 a_22250_772# VDD.t165 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X158 a_13406_352# en_4.t7 VSS.t70 VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X159 VDD.t8 en_0.t6 a_2496_772# VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X160 variable_delay_unit_2.in.t1 variable_delay_unit_1.in.t4 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X161 a_10458_772# variable_delay_unit_3.tristate_inverter_1.en.t6 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X162 variable_delay_unit_8.forward.t0 variable_delay_unit_8.in.t4 VSS.t97 VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X163 VSS.t88 variable_delay_unit_6.tristate_inverter_1.en.t6 a_20184_352# VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X164 variable_delay_unit_6.tristate_inverter_1.en.t1 en_6.t6 VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X165 VSS.t72 VDD.t169 a_25198_352# VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X166 variable_delay_unit_7.out variable_delay_unit_8.in.t5 a_22250_352# VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X167 variable_delay_unit_2.in.t0 variable_delay_unit_1.in.t5 VSS.t103 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X168 VSS.t124 variable_delay_unit_0.tristate_inverter_1.en.t6 a_2496_352# VSS.t123 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X169 VDD.t148 variable_delay_unit_7.tristate_inverter_1.en.t7 a_22250_772# VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X170 variable_delay_unit_6.tristate_inverter_1.en.t0 en_6.t7 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X171 a_10458_352# en_3.t6 VSS.t140 VSS.t139 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X172 VDD.t120 variable_delay_unit_0.tristate_inverter_1.en.t7 a_1614_772# VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X173 VDD.t133 en_3.t7 a_11340_772# VDD.t132 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X174 VSS.t136 en_7.t7 a_22250_352# VSS.t135 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X175 VDD.t71 VDD.t69 a_26080_772# VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X176 a_19302_772# variable_delay_unit_6.tristate_inverter_1.en.t7 VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X177 VSS.t115 en_0.t7 a_1614_352# VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X178 VSS.t84 variable_delay_unit_3.tristate_inverter_1.en.t7 a_11340_352# VSS.t83 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X179 VDD.t139 en_2.t7 a_8392_772# VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
R0 VDD.n448 VDD.n414 1689.71
R1 VDD.n419 VDD.n414 1689.71
R2 VDD.n412 VDD.n411 1689.71
R3 VDD.n451 VDD.n411 1689.71
R4 VDD.n388 VDD.n13 1689.71
R5 VDD.n388 VDD.n14 1689.71
R6 VDD.n20 VDD.n15 1689.71
R7 VDD.n384 VDD.n15 1689.71
R8 VDD.n360 VDD.n35 1689.71
R9 VDD.n360 VDD.n36 1689.71
R10 VDD.n42 VDD.n37 1689.71
R11 VDD.n356 VDD.n37 1689.71
R12 VDD.n332 VDD.n57 1689.71
R13 VDD.n332 VDD.n58 1689.71
R14 VDD.n64 VDD.n59 1689.71
R15 VDD.n328 VDD.n59 1689.71
R16 VDD.n304 VDD.n79 1689.71
R17 VDD.n304 VDD.n80 1689.71
R18 VDD.n86 VDD.n81 1689.71
R19 VDD.n300 VDD.n81 1689.71
R20 VDD.n276 VDD.n101 1689.71
R21 VDD.n276 VDD.n102 1689.71
R22 VDD.n108 VDD.n103 1689.71
R23 VDD.n272 VDD.n103 1689.71
R24 VDD.n248 VDD.n123 1689.71
R25 VDD.n248 VDD.n124 1689.71
R26 VDD.n130 VDD.n125 1689.71
R27 VDD.n244 VDD.n125 1689.71
R28 VDD.n220 VDD.n145 1689.71
R29 VDD.n220 VDD.n146 1689.71
R30 VDD.n152 VDD.n147 1689.71
R31 VDD.n216 VDD.n147 1689.71
R32 VDD.n184 VDD.n167 1689.71
R33 VDD.n184 VDD.n168 1689.71
R34 VDD.n174 VDD.n169 1689.71
R35 VDD.n180 VDD.n169 1689.71
R36 VDD.n198 VDD.n157 1307.92
R37 VDD.n194 VDD.n158 1307.92
R38 VDD.n234 VDD.n135 1307.92
R39 VDD.n230 VDD.n136 1307.92
R40 VDD.n262 VDD.n113 1307.92
R41 VDD.n258 VDD.n114 1307.92
R42 VDD.n290 VDD.n91 1307.92
R43 VDD.n286 VDD.n92 1307.92
R44 VDD.n318 VDD.n69 1307.92
R45 VDD.n314 VDD.n70 1307.92
R46 VDD.n346 VDD.n47 1307.92
R47 VDD.n342 VDD.n48 1307.92
R48 VDD.n374 VDD.n25 1307.92
R49 VDD.n370 VDD.n26 1307.92
R50 VDD.n402 VDD.n3 1307.92
R51 VDD.n398 VDD.n4 1307.92
R52 VDD.n431 VDD.n427 1307.92
R53 VDD.n424 VDD.n423 1307.92
R54 VDD.n204 VDD.t69 628.097
R55 VDD.n205 VDD.t72 622.766
R56 VDD.n208 VDD.t78 543.053
R57 VDD.n204 VDD.t75 523.774
R58 VDD.n450 VDD.n449 332.803
R59 VDD.n386 VDD.n385 332.803
R60 VDD.n358 VDD.n357 332.803
R61 VDD.n330 VDD.n329 332.803
R62 VDD.n302 VDD.n301 332.803
R63 VDD.n274 VDD.n273 332.803
R64 VDD.n246 VDD.n245 332.803
R65 VDD.n218 VDD.n217 332.803
R66 VDD.n182 VDD.n181 332.803
R67 VDD.n203 VDD.t166 304.647
R68 VDD.n203 VDD.t168 304.647
R69 VDD.n208 VDD.t167 221.72
R70 VDD.n209 VDD.n208 219.48
R71 VDD.n203 VDD.t169 202.44
R72 VDD.n447 VDD.n415 180.236
R73 VDD.n420 VDD.n415 180.236
R74 VDD.n453 VDD.n452 180.236
R75 VDD.n453 VDD.n407 180.236
R76 VDD.n389 VDD.n12 180.236
R77 VDD.n389 VDD.n8 180.236
R78 VDD.n383 VDD.n16 180.236
R79 VDD.n21 VDD.n16 180.236
R80 VDD.n361 VDD.n34 180.236
R81 VDD.n361 VDD.n30 180.236
R82 VDD.n355 VDD.n38 180.236
R83 VDD.n43 VDD.n38 180.236
R84 VDD.n333 VDD.n56 180.236
R85 VDD.n333 VDD.n52 180.236
R86 VDD.n327 VDD.n60 180.236
R87 VDD.n65 VDD.n60 180.236
R88 VDD.n305 VDD.n78 180.236
R89 VDD.n305 VDD.n74 180.236
R90 VDD.n299 VDD.n82 180.236
R91 VDD.n87 VDD.n82 180.236
R92 VDD.n277 VDD.n100 180.236
R93 VDD.n277 VDD.n96 180.236
R94 VDD.n271 VDD.n104 180.236
R95 VDD.n109 VDD.n104 180.236
R96 VDD.n249 VDD.n122 180.236
R97 VDD.n249 VDD.n118 180.236
R98 VDD.n243 VDD.n126 180.236
R99 VDD.n131 VDD.n126 180.236
R100 VDD.n221 VDD.n144 180.236
R101 VDD.n221 VDD.n140 180.236
R102 VDD.n215 VDD.n148 180.236
R103 VDD.n153 VDD.n148 180.236
R104 VDD.n185 VDD.n166 180.236
R105 VDD.n185 VDD.n162 180.236
R106 VDD.n179 VDD.n170 180.236
R107 VDD.n175 VDD.n170 180.236
R108 VDD.n197 VDD.n154 175.123
R109 VDD.n161 VDD.n160 175.123
R110 VDD.n233 VDD.n132 175.123
R111 VDD.n139 VDD.n138 175.123
R112 VDD.n261 VDD.n110 175.123
R113 VDD.n117 VDD.n116 175.123
R114 VDD.n289 VDD.n88 175.123
R115 VDD.n95 VDD.n94 175.123
R116 VDD.n317 VDD.n66 175.123
R117 VDD.n73 VDD.n72 175.123
R118 VDD.n345 VDD.n44 175.123
R119 VDD.n51 VDD.n50 175.123
R120 VDD.n373 VDD.n22 175.123
R121 VDD.n29 VDD.n28 175.123
R122 VDD.n401 VDD.n0 175.123
R123 VDD.n7 VDD.n6 175.123
R124 VDD.n434 VDD.n433 175.123
R125 VDD.n429 VDD.n421 175.123
R126 VDD VDD.n203 168.969
R127 VDD VDD.n205 166.147
R128 VDD.t130 VDD.n412 163.724
R129 VDD.n419 VDD.t44 163.724
R130 VDD.n20 VDD.t57 163.724
R131 VDD.t48 VDD.n14 163.724
R132 VDD.n42 VDD.t136 163.724
R133 VDD.t35 VDD.n36 163.724
R134 VDD.n64 VDD.t65 163.724
R135 VDD.t149 VDD.n58 163.724
R136 VDD.n86 VDD.t18 163.724
R137 VDD.t40 VDD.n80 163.724
R138 VDD.n108 VDD.t67 163.724
R139 VDD.t12 VDD.n102 163.724
R140 VDD.n130 VDD.t90 163.724
R141 VDD.t22 VDD.n124 163.724
R142 VDD.n152 VDD.t125 163.724
R143 VDD.t123 VDD.n146 163.724
R144 VDD.n174 VDD.t70 163.724
R145 VDD.t121 VDD.n168 163.724
R146 VDD.n195 VDD.t162 160.923
R147 VDD.t79 VDD.n196 160.923
R148 VDD.n231 VDD.t86 160.923
R149 VDD.t38 VDD.n232 160.923
R150 VDD.n259 VDD.t30 160.923
R151 VDD.t140 VDD.n260 160.923
R152 VDD.n287 VDD.t25 160.923
R153 VDD.t0 VDD.n288 160.923
R154 VDD.n315 VDD.t59 160.923
R155 VDD.t92 VDD.n316 160.923
R156 VDD.n343 VDD.t142 160.923
R157 VDD.t61 VDD.n344 160.923
R158 VDD.n371 VDD.t42 160.923
R159 VDD.t160 VDD.n372 160.923
R160 VDD.n399 VDD.t108 160.923
R161 VDD.t152 VDD.n400 160.923
R162 VDD.n430 VDD.t4 160.923
R163 VDD.t88 VDD.n432 160.923
R164 VDD.n450 VDD.t151 145.224
R165 VDD.n449 VDD.t9 145.224
R166 VDD.n385 VDD.t114 145.224
R167 VDD.t146 VDD.n386 145.224
R168 VDD.n357 VDD.t145 145.224
R169 VDD.t83 VDD.n358 145.224
R170 VDD.n329 VDD.t98 145.224
R171 VDD.t144 VDD.n330 145.224
R172 VDD.n301 VDD.t6 145.224
R173 VDD.t24 VDD.n302 145.224
R174 VDD.n273 VDD.t37 145.224
R175 VDD.t29 VDD.n274 145.224
R176 VDD.n245 VDD.t105 145.224
R177 VDD.t164 VDD.n246 145.224
R178 VDD.n217 VDD.t50 145.224
R179 VDD.t165 VDD.n218 145.224
R180 VDD.n181 VDD.t34 145.224
R181 VDD.t129 VDD.n182 145.224
R182 VDD.n199 VDD.n156 139.512
R183 VDD.n199 VDD.n154 139.512
R184 VDD.n193 VDD.n159 139.512
R185 VDD.n161 VDD.n159 139.512
R186 VDD.n235 VDD.n134 139.512
R187 VDD.n235 VDD.n132 139.512
R188 VDD.n229 VDD.n137 139.512
R189 VDD.n139 VDD.n137 139.512
R190 VDD.n263 VDD.n112 139.512
R191 VDD.n263 VDD.n110 139.512
R192 VDD.n257 VDD.n115 139.512
R193 VDD.n117 VDD.n115 139.512
R194 VDD.n291 VDD.n90 139.512
R195 VDD.n291 VDD.n88 139.512
R196 VDD.n285 VDD.n93 139.512
R197 VDD.n95 VDD.n93 139.512
R198 VDD.n319 VDD.n68 139.512
R199 VDD.n319 VDD.n66 139.512
R200 VDD.n313 VDD.n71 139.512
R201 VDD.n73 VDD.n71 139.512
R202 VDD.n347 VDD.n46 139.512
R203 VDD.n347 VDD.n44 139.512
R204 VDD.n341 VDD.n49 139.512
R205 VDD.n51 VDD.n49 139.512
R206 VDD.n375 VDD.n24 139.512
R207 VDD.n375 VDD.n22 139.512
R208 VDD.n369 VDD.n27 139.512
R209 VDD.n29 VDD.n27 139.512
R210 VDD.n403 VDD.n2 139.512
R211 VDD.n403 VDD.n0 139.512
R212 VDD.n397 VDD.n5 139.512
R213 VDD.n7 VDD.n5 139.512
R214 VDD.n435 VDD.n425 139.512
R215 VDD.n435 VDD.n434 139.512
R216 VDD.n440 VDD.n439 139.512
R217 VDD.n440 VDD.n421 139.512
R218 VDD.n196 VDD.n195 119.861
R219 VDD.n232 VDD.n231 119.861
R220 VDD.n260 VDD.n259 119.861
R221 VDD.n288 VDD.n287 119.861
R222 VDD.n316 VDD.n315 119.861
R223 VDD.n344 VDD.n343 119.861
R224 VDD.n372 VDD.n371 119.861
R225 VDD.n400 VDD.n399 119.861
R226 VDD.n432 VDD.n430 119.861
R227 VDD.t110 VDD.t130 88.7478
R228 VDD.t151 VDD.t7 88.7478
R229 VDD.t103 VDD.t9 88.7478
R230 VDD.t44 VDD.t119 88.7478
R231 VDD.t57 VDD.t84 88.7478
R232 VDD.t53 VDD.t114 88.7478
R233 VDD.t32 VDD.t146 88.7478
R234 VDD.t156 VDD.t48 88.7478
R235 VDD.t136 VDD.t158 88.7478
R236 VDD.t138 VDD.t145 88.7478
R237 VDD.t154 VDD.t83 88.7478
R238 VDD.t101 VDD.t35 88.7478
R239 VDD.t65 VDD.t63 88.7478
R240 VDD.t132 VDD.t98 88.7478
R241 VDD.t106 VDD.t144 88.7478
R242 VDD.t115 VDD.t149 88.7478
R243 VDD.t18 VDD.t46 88.7478
R244 VDD.t20 VDD.t6 88.7478
R245 VDD.t96 VDD.t24 88.7478
R246 VDD.t81 VDD.t40 88.7478
R247 VDD.t67 VDD.t2 88.7478
R248 VDD.t55 VDD.t37 88.7478
R249 VDD.t99 VDD.t29 88.7478
R250 VDD.t51 VDD.t12 88.7478
R251 VDD.t90 VDD.t27 88.7478
R252 VDD.t16 VDD.t105 88.7478
R253 VDD.t117 VDD.t164 88.7478
R254 VDD.t134 VDD.t22 88.7478
R255 VDD.t125 VDD.t112 88.7478
R256 VDD.t127 VDD.t50 88.7478
R257 VDD.t94 VDD.t165 88.7478
R258 VDD.t147 VDD.t123 88.7478
R259 VDD.t70 VDD.t76 88.7478
R260 VDD.t73 VDD.t34 88.7478
R261 VDD.t10 VDD.t129 88.7478
R262 VDD.t14 VDD.t121 88.7478
R263 VDD.n201 VDD.t80 84.7934
R264 VDD.n191 VDD.t163 84.7934
R265 VDD.n237 VDD.t39 84.7934
R266 VDD.n227 VDD.t87 84.7934
R267 VDD.n265 VDD.t141 84.7934
R268 VDD.n255 VDD.t31 84.7934
R269 VDD.n293 VDD.t1 84.7934
R270 VDD.n283 VDD.t26 84.7934
R271 VDD.n321 VDD.t93 84.7934
R272 VDD.n311 VDD.t60 84.7934
R273 VDD.n349 VDD.t62 84.7934
R274 VDD.n339 VDD.t143 84.7934
R275 VDD.n377 VDD.t161 84.7934
R276 VDD.n367 VDD.t43 84.7934
R277 VDD.n405 VDD.t153 84.7934
R278 VDD.n395 VDD.t109 84.7934
R279 VDD.n426 VDD.t89 84.7934
R280 VDD.n422 VDD.t5 84.7934
R281 VDD.n417 VDD.n416 84.7744
R282 VDD.n409 VDD.n408 84.7744
R283 VDD.n10 VDD.n9 84.7744
R284 VDD.n18 VDD.n17 84.7744
R285 VDD.n32 VDD.n31 84.7744
R286 VDD.n40 VDD.n39 84.7744
R287 VDD.n54 VDD.n53 84.7744
R288 VDD.n62 VDD.n61 84.7744
R289 VDD.n76 VDD.n75 84.7744
R290 VDD.n84 VDD.n83 84.7744
R291 VDD.n98 VDD.n97 84.7744
R292 VDD.n106 VDD.n105 84.7744
R293 VDD.n120 VDD.n119 84.7744
R294 VDD.n128 VDD.n127 84.7744
R295 VDD.n142 VDD.n141 84.7744
R296 VDD.n150 VDD.n149 84.7744
R297 VDD.n164 VDD.n163 84.7744
R298 VDD.n172 VDD.n171 84.7744
R299 VDD.n417 VDD.t45 83.8097
R300 VDD.n409 VDD.t131 83.8097
R301 VDD.n10 VDD.t49 83.8097
R302 VDD.n18 VDD.t58 83.8097
R303 VDD.n32 VDD.t36 83.8097
R304 VDD.n40 VDD.t137 83.8097
R305 VDD.n54 VDD.t150 83.8097
R306 VDD.n62 VDD.t66 83.8097
R307 VDD.n76 VDD.t41 83.8097
R308 VDD.n84 VDD.t19 83.8097
R309 VDD.n98 VDD.t13 83.8097
R310 VDD.n106 VDD.t68 83.8097
R311 VDD.n120 VDD.t23 83.8097
R312 VDD.n128 VDD.t91 83.8097
R313 VDD.n142 VDD.t124 83.8097
R314 VDD.n150 VDD.t126 83.8097
R315 VDD.n164 VDD.t122 83.8097
R316 VDD.n172 VDD.t71 83.8097
R317 VDD.n199 VDD.n198 46.2505
R318 VDD.n159 VDD.n158 46.2505
R319 VDD.n235 VDD.n234 46.2505
R320 VDD.n137 VDD.n136 46.2505
R321 VDD.n263 VDD.n262 46.2505
R322 VDD.n115 VDD.n114 46.2505
R323 VDD.n291 VDD.n290 46.2505
R324 VDD.n93 VDD.n92 46.2505
R325 VDD.n319 VDD.n318 46.2505
R326 VDD.n71 VDD.n70 46.2505
R327 VDD.n347 VDD.n346 46.2505
R328 VDD.n49 VDD.n48 46.2505
R329 VDD.n375 VDD.n374 46.2505
R330 VDD.n27 VDD.n26 46.2505
R331 VDD.n403 VDD.n402 46.2505
R332 VDD.n5 VDD.n4 46.2505
R333 VDD.n435 VDD.n427 46.2505
R334 VDD.n440 VDD.n423 46.2505
R335 VDD.n413 VDD.t110 44.3742
R336 VDD.t7 VDD.n413 44.3742
R337 VDD.n418 VDD.t103 44.3742
R338 VDD.t119 VDD.n418 44.3742
R339 VDD.t84 VDD.n19 44.3742
R340 VDD.n19 VDD.t53 44.3742
R341 VDD.n387 VDD.t32 44.3742
R342 VDD.n387 VDD.t156 44.3742
R343 VDD.t158 VDD.n41 44.3742
R344 VDD.n41 VDD.t138 44.3742
R345 VDD.n359 VDD.t154 44.3742
R346 VDD.n359 VDD.t101 44.3742
R347 VDD.t63 VDD.n63 44.3742
R348 VDD.n63 VDD.t132 44.3742
R349 VDD.n331 VDD.t106 44.3742
R350 VDD.n331 VDD.t115 44.3742
R351 VDD.t46 VDD.n85 44.3742
R352 VDD.n85 VDD.t20 44.3742
R353 VDD.n303 VDD.t96 44.3742
R354 VDD.n303 VDD.t81 44.3742
R355 VDD.t2 VDD.n107 44.3742
R356 VDD.n107 VDD.t55 44.3742
R357 VDD.n275 VDD.t99 44.3742
R358 VDD.n275 VDD.t51 44.3742
R359 VDD.t27 VDD.n129 44.3742
R360 VDD.n129 VDD.t16 44.3742
R361 VDD.n247 VDD.t117 44.3742
R362 VDD.n247 VDD.t134 44.3742
R363 VDD.t112 VDD.n151 44.3742
R364 VDD.n151 VDD.t127 44.3742
R365 VDD.n219 VDD.t94 44.3742
R366 VDD.n219 VDD.t147 44.3742
R367 VDD.t76 VDD.n173 44.3742
R368 VDD.n173 VDD.t73 44.3742
R369 VDD.n183 VDD.t10 44.3742
R370 VDD.n183 VDD.t14 44.3742
R371 VDD.n198 VDD.n197 39.3924
R372 VDD.n160 VDD.n158 39.3924
R373 VDD.n234 VDD.n233 39.3924
R374 VDD.n138 VDD.n136 39.3924
R375 VDD.n262 VDD.n261 39.3924
R376 VDD.n116 VDD.n114 39.3924
R377 VDD.n290 VDD.n289 39.3924
R378 VDD.n94 VDD.n92 39.3924
R379 VDD.n318 VDD.n317 39.3924
R380 VDD.n72 VDD.n70 39.3924
R381 VDD.n346 VDD.n345 39.3924
R382 VDD.n50 VDD.n48 39.3924
R383 VDD.n374 VDD.n373 39.3924
R384 VDD.n28 VDD.n26 39.3924
R385 VDD.n402 VDD.n401 39.3924
R386 VDD.n6 VDD.n4 39.3924
R387 VDD.n433 VDD.n427 39.3924
R388 VDD.n429 VDD.n423 39.3924
R389 VDD.n415 VDD.n414 23.1255
R390 VDD.n418 VDD.n414 23.1255
R391 VDD.n453 VDD.n411 23.1255
R392 VDD.n413 VDD.n411 23.1255
R393 VDD.n389 VDD.n388 23.1255
R394 VDD.n388 VDD.n387 23.1255
R395 VDD.n16 VDD.n15 23.1255
R396 VDD.n19 VDD.n15 23.1255
R397 VDD.n361 VDD.n360 23.1255
R398 VDD.n360 VDD.n359 23.1255
R399 VDD.n38 VDD.n37 23.1255
R400 VDD.n41 VDD.n37 23.1255
R401 VDD.n333 VDD.n332 23.1255
R402 VDD.n332 VDD.n331 23.1255
R403 VDD.n60 VDD.n59 23.1255
R404 VDD.n63 VDD.n59 23.1255
R405 VDD.n305 VDD.n304 23.1255
R406 VDD.n304 VDD.n303 23.1255
R407 VDD.n82 VDD.n81 23.1255
R408 VDD.n85 VDD.n81 23.1255
R409 VDD.n277 VDD.n276 23.1255
R410 VDD.n276 VDD.n275 23.1255
R411 VDD.n104 VDD.n103 23.1255
R412 VDD.n107 VDD.n103 23.1255
R413 VDD.n249 VDD.n248 23.1255
R414 VDD.n248 VDD.n247 23.1255
R415 VDD.n126 VDD.n125 23.1255
R416 VDD.n129 VDD.n125 23.1255
R417 VDD.n221 VDD.n220 23.1255
R418 VDD.n220 VDD.n219 23.1255
R419 VDD.n148 VDD.n147 23.1255
R420 VDD.n151 VDD.n147 23.1255
R421 VDD.n185 VDD.n184 23.1255
R422 VDD.n184 VDD.n183 23.1255
R423 VDD.n170 VDD.n169 23.1255
R424 VDD.n173 VDD.n169 23.1255
R425 VDD.n157 VDD.n156 20.5561
R426 VDD.n196 VDD.n157 20.5561
R427 VDD.n194 VDD.n193 20.5561
R428 VDD.n195 VDD.n194 20.5561
R429 VDD.n135 VDD.n134 20.5561
R430 VDD.n232 VDD.n135 20.5561
R431 VDD.n230 VDD.n229 20.5561
R432 VDD.n231 VDD.n230 20.5561
R433 VDD.n113 VDD.n112 20.5561
R434 VDD.n260 VDD.n113 20.5561
R435 VDD.n258 VDD.n257 20.5561
R436 VDD.n259 VDD.n258 20.5561
R437 VDD.n91 VDD.n90 20.5561
R438 VDD.n288 VDD.n91 20.5561
R439 VDD.n286 VDD.n285 20.5561
R440 VDD.n287 VDD.n286 20.5561
R441 VDD.n69 VDD.n68 20.5561
R442 VDD.n316 VDD.n69 20.5561
R443 VDD.n314 VDD.n313 20.5561
R444 VDD.n315 VDD.n314 20.5561
R445 VDD.n47 VDD.n46 20.5561
R446 VDD.n344 VDD.n47 20.5561
R447 VDD.n342 VDD.n341 20.5561
R448 VDD.n343 VDD.n342 20.5561
R449 VDD.n25 VDD.n24 20.5561
R450 VDD.n372 VDD.n25 20.5561
R451 VDD.n370 VDD.n369 20.5561
R452 VDD.n371 VDD.n370 20.5561
R453 VDD.n3 VDD.n2 20.5561
R454 VDD.n400 VDD.n3 20.5561
R455 VDD.n398 VDD.n397 20.5561
R456 VDD.n399 VDD.n398 20.5561
R457 VDD.n431 VDD.n425 20.5561
R458 VDD.n432 VDD.n431 20.5561
R459 VDD.n439 VDD.n424 20.5561
R460 VDD.n430 VDD.n424 20.5561
R461 VDD.n420 VDD.n419 18.5005
R462 VDD.n448 VDD.n447 18.5005
R463 VDD.n449 VDD.n448 18.5005
R464 VDD.n452 VDD.n451 18.5005
R465 VDD.n451 VDD.n450 18.5005
R466 VDD.n412 VDD.n407 18.5005
R467 VDD.n14 VDD.n8 18.5005
R468 VDD.n13 VDD.n12 18.5005
R469 VDD.n386 VDD.n13 18.5005
R470 VDD.n384 VDD.n383 18.5005
R471 VDD.n385 VDD.n384 18.5005
R472 VDD.n21 VDD.n20 18.5005
R473 VDD.n36 VDD.n30 18.5005
R474 VDD.n35 VDD.n34 18.5005
R475 VDD.n358 VDD.n35 18.5005
R476 VDD.n356 VDD.n355 18.5005
R477 VDD.n357 VDD.n356 18.5005
R478 VDD.n43 VDD.n42 18.5005
R479 VDD.n58 VDD.n52 18.5005
R480 VDD.n57 VDD.n56 18.5005
R481 VDD.n330 VDD.n57 18.5005
R482 VDD.n328 VDD.n327 18.5005
R483 VDD.n329 VDD.n328 18.5005
R484 VDD.n65 VDD.n64 18.5005
R485 VDD.n80 VDD.n74 18.5005
R486 VDD.n79 VDD.n78 18.5005
R487 VDD.n302 VDD.n79 18.5005
R488 VDD.n300 VDD.n299 18.5005
R489 VDD.n301 VDD.n300 18.5005
R490 VDD.n87 VDD.n86 18.5005
R491 VDD.n102 VDD.n96 18.5005
R492 VDD.n101 VDD.n100 18.5005
R493 VDD.n274 VDD.n101 18.5005
R494 VDD.n272 VDD.n271 18.5005
R495 VDD.n273 VDD.n272 18.5005
R496 VDD.n109 VDD.n108 18.5005
R497 VDD.n124 VDD.n118 18.5005
R498 VDD.n123 VDD.n122 18.5005
R499 VDD.n246 VDD.n123 18.5005
R500 VDD.n244 VDD.n243 18.5005
R501 VDD.n245 VDD.n244 18.5005
R502 VDD.n131 VDD.n130 18.5005
R503 VDD.n146 VDD.n140 18.5005
R504 VDD.n145 VDD.n144 18.5005
R505 VDD.n218 VDD.n145 18.5005
R506 VDD.n216 VDD.n215 18.5005
R507 VDD.n217 VDD.n216 18.5005
R508 VDD.n153 VDD.n152 18.5005
R509 VDD.n168 VDD.n162 18.5005
R510 VDD.n167 VDD.n166 18.5005
R511 VDD.n182 VDD.n167 18.5005
R512 VDD.n180 VDD.n179 18.5005
R513 VDD.n181 VDD.n180 18.5005
R514 VDD.n175 VDD.n174 18.5005
R515 VDD.n416 VDD.t104 9.52217
R516 VDD.n416 VDD.t120 9.52217
R517 VDD.n408 VDD.t111 9.52217
R518 VDD.n408 VDD.t8 9.52217
R519 VDD.n9 VDD.t33 9.52217
R520 VDD.n9 VDD.t157 9.52217
R521 VDD.n17 VDD.t85 9.52217
R522 VDD.n17 VDD.t54 9.52217
R523 VDD.n31 VDD.t155 9.52217
R524 VDD.n31 VDD.t102 9.52217
R525 VDD.n39 VDD.t159 9.52217
R526 VDD.n39 VDD.t139 9.52217
R527 VDD.n53 VDD.t107 9.52217
R528 VDD.n53 VDD.t116 9.52217
R529 VDD.n61 VDD.t64 9.52217
R530 VDD.n61 VDD.t133 9.52217
R531 VDD.n75 VDD.t97 9.52217
R532 VDD.n75 VDD.t82 9.52217
R533 VDD.n83 VDD.t47 9.52217
R534 VDD.n83 VDD.t21 9.52217
R535 VDD.n97 VDD.t100 9.52217
R536 VDD.n97 VDD.t52 9.52217
R537 VDD.n105 VDD.t3 9.52217
R538 VDD.n105 VDD.t56 9.52217
R539 VDD.n119 VDD.t118 9.52217
R540 VDD.n119 VDD.t135 9.52217
R541 VDD.n127 VDD.t28 9.52217
R542 VDD.n127 VDD.t17 9.52217
R543 VDD.n141 VDD.t95 9.52217
R544 VDD.n141 VDD.t148 9.52217
R545 VDD.n149 VDD.t113 9.52217
R546 VDD.n149 VDD.t128 9.52217
R547 VDD.n163 VDD.t11 9.52217
R548 VDD.n163 VDD.t15 9.52217
R549 VDD.n171 VDD.t77 9.52217
R550 VDD.n171 VDD.t74 9.52217
R551 VDD.n160 VDD.t162 5.4667
R552 VDD.n197 VDD.t79 5.4667
R553 VDD.n138 VDD.t86 5.4667
R554 VDD.n233 VDD.t38 5.4667
R555 VDD.n116 VDD.t30 5.4667
R556 VDD.n261 VDD.t140 5.4667
R557 VDD.n94 VDD.t25 5.4667
R558 VDD.n289 VDD.t0 5.4667
R559 VDD.n72 VDD.t59 5.4667
R560 VDD.n317 VDD.t92 5.4667
R561 VDD.n50 VDD.t142 5.4667
R562 VDD.n345 VDD.t61 5.4667
R563 VDD.n28 VDD.t42 5.4667
R564 VDD.n373 VDD.t160 5.4667
R565 VDD.n6 VDD.t108 5.4667
R566 VDD.n401 VDD.t152 5.4667
R567 VDD.t4 VDD.n429 5.4667
R568 VDD.n433 VDD.t88 5.4667
R569 VDD.n210 VDD.n209 4.5005
R570 VDD.n207 VDD.n206 3.26479
R571 VDD.n190 VDD.n159 2.3255
R572 VDD.n200 VDD.n199 2.3255
R573 VDD.n226 VDD.n137 2.3255
R574 VDD.n236 VDD.n235 2.3255
R575 VDD.n254 VDD.n115 2.3255
R576 VDD.n264 VDD.n263 2.3255
R577 VDD.n282 VDD.n93 2.3255
R578 VDD.n292 VDD.n291 2.3255
R579 VDD.n310 VDD.n71 2.3255
R580 VDD.n320 VDD.n319 2.3255
R581 VDD.n338 VDD.n49 2.3255
R582 VDD.n348 VDD.n347 2.3255
R583 VDD.n366 VDD.n27 2.3255
R584 VDD.n376 VDD.n375 2.3255
R585 VDD.n394 VDD.n5 2.3255
R586 VDD.n404 VDD.n403 2.3255
R587 VDD.n441 VDD.n440 2.3255
R588 VDD.n436 VDD.n435 2.3255
R589 VDD.n193 VDD.n192 2.04321
R590 VDD.n202 VDD.n154 2.04321
R591 VDD.n156 VDD.n155 2.04321
R592 VDD.n189 VDD.n161 2.04321
R593 VDD.n229 VDD.n228 2.04321
R594 VDD.n238 VDD.n132 2.04321
R595 VDD.n134 VDD.n133 2.04321
R596 VDD.n225 VDD.n139 2.04321
R597 VDD.n257 VDD.n256 2.04321
R598 VDD.n266 VDD.n110 2.04321
R599 VDD.n112 VDD.n111 2.04321
R600 VDD.n253 VDD.n117 2.04321
R601 VDD.n285 VDD.n284 2.04321
R602 VDD.n294 VDD.n88 2.04321
R603 VDD.n90 VDD.n89 2.04321
R604 VDD.n281 VDD.n95 2.04321
R605 VDD.n313 VDD.n312 2.04321
R606 VDD.n322 VDD.n66 2.04321
R607 VDD.n68 VDD.n67 2.04321
R608 VDD.n309 VDD.n73 2.04321
R609 VDD.n341 VDD.n340 2.04321
R610 VDD.n350 VDD.n44 2.04321
R611 VDD.n46 VDD.n45 2.04321
R612 VDD.n337 VDD.n51 2.04321
R613 VDD.n369 VDD.n368 2.04321
R614 VDD.n378 VDD.n22 2.04321
R615 VDD.n24 VDD.n23 2.04321
R616 VDD.n365 VDD.n29 2.04321
R617 VDD.n397 VDD.n396 2.04321
R618 VDD.n406 VDD.n0 2.04321
R619 VDD.n2 VDD.n1 2.04321
R620 VDD.n393 VDD.n7 2.04321
R621 VDD.n439 VDD.n438 2.04321
R622 VDD.n434 VDD.n428 2.04321
R623 VDD.n437 VDD.n425 2.04321
R624 VDD.n442 VDD.n421 2.04321
R625 VDD VDD.n175 1.97234
R626 VDD.n452 VDD.n410 1.96583
R627 VDD.n443 VDD.n420 1.96583
R628 VDD.n447 VDD.n446 1.96583
R629 VDD.n456 VDD.n407 1.96583
R630 VDD.n383 VDD.n382 1.96583
R631 VDD.n392 VDD.n8 1.96583
R632 VDD.n12 VDD.n11 1.96583
R633 VDD.n379 VDD.n21 1.96583
R634 VDD.n355 VDD.n354 1.96583
R635 VDD.n364 VDD.n30 1.96583
R636 VDD.n34 VDD.n33 1.96583
R637 VDD.n351 VDD.n43 1.96583
R638 VDD.n327 VDD.n326 1.96583
R639 VDD.n336 VDD.n52 1.96583
R640 VDD.n56 VDD.n55 1.96583
R641 VDD.n323 VDD.n65 1.96583
R642 VDD.n299 VDD.n298 1.96583
R643 VDD.n308 VDD.n74 1.96583
R644 VDD.n78 VDD.n77 1.96583
R645 VDD.n295 VDD.n87 1.96583
R646 VDD.n271 VDD.n270 1.96583
R647 VDD.n280 VDD.n96 1.96583
R648 VDD.n100 VDD.n99 1.96583
R649 VDD.n267 VDD.n109 1.96583
R650 VDD.n243 VDD.n242 1.96583
R651 VDD.n252 VDD.n118 1.96583
R652 VDD.n122 VDD.n121 1.96583
R653 VDD.n239 VDD.n131 1.96583
R654 VDD.n215 VDD.n214 1.96583
R655 VDD.n224 VDD.n140 1.96583
R656 VDD.n144 VDD.n143 1.96583
R657 VDD.n211 VDD.n153 1.96583
R658 VDD.n179 VDD.n178 1.96583
R659 VDD.n188 VDD.n162 1.96583
R660 VDD.n166 VDD.n165 1.96583
R661 VDD.n206 VDD 1.40175
R662 VDD.n177 VDD.n170 1.32907
R663 VDD.n186 VDD.n185 1.32907
R664 VDD.n213 VDD.n148 1.32907
R665 VDD.n222 VDD.n221 1.32907
R666 VDD.n241 VDD.n126 1.32907
R667 VDD.n250 VDD.n249 1.32907
R668 VDD.n269 VDD.n104 1.32907
R669 VDD.n278 VDD.n277 1.32907
R670 VDD.n297 VDD.n82 1.32907
R671 VDD.n306 VDD.n305 1.32907
R672 VDD.n325 VDD.n60 1.32907
R673 VDD.n334 VDD.n333 1.32907
R674 VDD.n353 VDD.n38 1.32907
R675 VDD.n362 VDD.n361 1.32907
R676 VDD.n381 VDD.n16 1.32907
R677 VDD.n390 VDD.n389 1.32907
R678 VDD.n454 VDD.n453 1.32907
R679 VDD.n445 VDD.n415 1.32907
R680 VDD.n444 VDD.n417 1.21789
R681 VDD.n455 VDD.n409 1.21789
R682 VDD.n391 VDD.n10 1.21789
R683 VDD.n380 VDD.n18 1.21789
R684 VDD.n363 VDD.n32 1.21789
R685 VDD.n352 VDD.n40 1.21789
R686 VDD.n335 VDD.n54 1.21789
R687 VDD.n324 VDD.n62 1.21789
R688 VDD.n307 VDD.n76 1.21789
R689 VDD.n296 VDD.n84 1.21789
R690 VDD.n279 VDD.n98 1.21789
R691 VDD.n268 VDD.n106 1.21789
R692 VDD.n251 VDD.n120 1.21789
R693 VDD.n240 VDD.n128 1.21789
R694 VDD.n223 VDD.n142 1.21789
R695 VDD.n212 VDD.n150 1.21789
R696 VDD.n187 VDD.n164 1.21789
R697 VDD.n176 VDD.n172 1.21789
R698 VDD.n205 VDD.n204 1.09595
R699 VDD.n209 VDD.n207 0.784429
R700 VDD VDD.n238 0.568208
R701 VDD VDD.n266 0.568208
R702 VDD VDD.n294 0.568208
R703 VDD VDD.n322 0.568208
R704 VDD VDD.n350 0.568208
R705 VDD VDD.n378 0.568208
R706 VDD VDD.n406 0.568208
R707 VDD.n428 VDD 0.492688
R708 VDD.n206 VDD 0.443357
R709 VDD.n189 VDD 0.432792
R710 VDD.n225 VDD 0.432792
R711 VDD.n253 VDD 0.432792
R712 VDD.n281 VDD 0.432792
R713 VDD.n309 VDD 0.432792
R714 VDD.n337 VDD 0.432792
R715 VDD.n365 VDD 0.432792
R716 VDD.n393 VDD 0.432792
R717 VDD VDD.n442 0.432792
R718 VDD.n178 VDD.n165 0.430188
R719 VDD.n214 VDD.n143 0.430188
R720 VDD.n242 VDD.n121 0.430188
R721 VDD.n270 VDD.n99 0.430188
R722 VDD.n298 VDD.n77 0.430188
R723 VDD.n326 VDD.n55 0.430188
R724 VDD.n354 VDD.n33 0.430188
R725 VDD.n382 VDD.n11 0.430188
R726 VDD.n446 VDD.n410 0.430188
R727 VDD VDD.n210 0.393729
R728 VDD.n178 VDD.n177 0.359875
R729 VDD.n186 VDD.n165 0.359875
R730 VDD.n214 VDD.n213 0.359875
R731 VDD.n222 VDD.n143 0.359875
R732 VDD.n242 VDD.n241 0.359875
R733 VDD.n250 VDD.n121 0.359875
R734 VDD.n270 VDD.n269 0.359875
R735 VDD.n278 VDD.n99 0.359875
R736 VDD.n298 VDD.n297 0.359875
R737 VDD.n306 VDD.n77 0.359875
R738 VDD.n326 VDD.n325 0.359875
R739 VDD.n334 VDD.n55 0.359875
R740 VDD.n354 VDD.n353 0.359875
R741 VDD.n362 VDD.n33 0.359875
R742 VDD.n382 VDD.n381 0.359875
R743 VDD.n390 VDD.n11 0.359875
R744 VDD.n454 VDD.n410 0.359875
R745 VDD.n446 VDD.n445 0.359875
R746 VDD.n177 VDD.n176 0.229667
R747 VDD.n187 VDD.n186 0.229667
R748 VDD.n213 VDD.n212 0.229667
R749 VDD.n223 VDD.n222 0.229667
R750 VDD.n241 VDD.n240 0.229667
R751 VDD.n251 VDD.n250 0.229667
R752 VDD.n269 VDD.n268 0.229667
R753 VDD.n279 VDD.n278 0.229667
R754 VDD.n297 VDD.n296 0.229667
R755 VDD.n307 VDD.n306 0.229667
R756 VDD.n325 VDD.n324 0.229667
R757 VDD.n335 VDD.n334 0.229667
R758 VDD.n353 VDD.n352 0.229667
R759 VDD.n363 VDD.n362 0.229667
R760 VDD.n381 VDD.n380 0.229667
R761 VDD.n391 VDD.n390 0.229667
R762 VDD.n455 VDD.n454 0.229667
R763 VDD.n445 VDD.n444 0.229667
R764 VDD.n190 VDD.n189 0.189302
R765 VDD.n200 VDD.n155 0.189302
R766 VDD.n226 VDD.n225 0.189302
R767 VDD.n236 VDD.n133 0.189302
R768 VDD.n254 VDD.n253 0.189302
R769 VDD.n264 VDD.n111 0.189302
R770 VDD.n282 VDD.n281 0.189302
R771 VDD.n292 VDD.n89 0.189302
R772 VDD.n310 VDD.n309 0.189302
R773 VDD.n320 VDD.n67 0.189302
R774 VDD.n338 VDD.n337 0.189302
R775 VDD.n348 VDD.n45 0.189302
R776 VDD.n366 VDD.n365 0.189302
R777 VDD.n376 VDD.n23 0.189302
R778 VDD.n394 VDD.n393 0.189302
R779 VDD.n404 VDD.n1 0.189302
R780 VDD.n442 VDD.n441 0.189302
R781 VDD.n437 VDD.n436 0.189302
R782 VDD.n210 VDD.n202 0.174979
R783 VDD.n192 VDD.n155 0.141125
R784 VDD.n228 VDD.n133 0.141125
R785 VDD.n256 VDD.n111 0.141125
R786 VDD.n284 VDD.n89 0.141125
R787 VDD.n312 VDD.n67 0.141125
R788 VDD.n340 VDD.n45 0.141125
R789 VDD.n368 VDD.n23 0.141125
R790 VDD.n396 VDD.n1 0.141125
R791 VDD.n438 VDD.n437 0.141125
R792 VDD.n192 VDD.n191 0.13201
R793 VDD.n202 VDD.n201 0.13201
R794 VDD.n228 VDD.n227 0.13201
R795 VDD.n238 VDD.n237 0.13201
R796 VDD.n256 VDD.n255 0.13201
R797 VDD.n266 VDD.n265 0.13201
R798 VDD.n284 VDD.n283 0.13201
R799 VDD.n294 VDD.n293 0.13201
R800 VDD.n312 VDD.n311 0.13201
R801 VDD.n322 VDD.n321 0.13201
R802 VDD.n340 VDD.n339 0.13201
R803 VDD.n350 VDD.n349 0.13201
R804 VDD.n368 VDD.n367 0.13201
R805 VDD.n378 VDD.n377 0.13201
R806 VDD.n396 VDD.n395 0.13201
R807 VDD.n406 VDD.n405 0.13201
R808 VDD.n438 VDD.n422 0.13201
R809 VDD.n428 VDD.n426 0.13201
R810 VDD.n188 VDD.n187 0.130708
R811 VDD.n224 VDD.n223 0.130708
R812 VDD.n252 VDD.n251 0.130708
R813 VDD.n280 VDD.n279 0.130708
R814 VDD.n308 VDD.n307 0.130708
R815 VDD.n336 VDD.n335 0.130708
R816 VDD.n364 VDD.n363 0.130708
R817 VDD.n392 VDD.n391 0.130708
R818 VDD.n444 VDD.n443 0.130708
R819 VDD.n176 VDD 0.124198
R820 VDD.n212 VDD 0.124198
R821 VDD.n240 VDD 0.124198
R822 VDD.n268 VDD 0.124198
R823 VDD.n296 VDD 0.124198
R824 VDD.n324 VDD 0.124198
R825 VDD.n352 VDD 0.124198
R826 VDD.n380 VDD 0.124198
R827 VDD VDD.n455 0.124198
R828 VDD VDD.n188 0.0695104
R829 VDD.n211 VDD 0.0695104
R830 VDD VDD.n224 0.0695104
R831 VDD.n239 VDD 0.0695104
R832 VDD VDD.n252 0.0695104
R833 VDD.n267 VDD 0.0695104
R834 VDD VDD.n280 0.0695104
R835 VDD.n295 VDD 0.0695104
R836 VDD VDD.n308 0.0695104
R837 VDD.n323 VDD 0.0695104
R838 VDD VDD.n336 0.0695104
R839 VDD.n351 VDD 0.0695104
R840 VDD VDD.n364 0.0695104
R841 VDD.n379 VDD 0.0695104
R842 VDD VDD.n392 0.0695104
R843 VDD VDD.n456 0.0695104
R844 VDD.n443 VDD 0.0695104
R845 VDD.n207 VDD 0.063
R846 VDD.n191 VDD.n190 0.0577917
R847 VDD.n201 VDD.n200 0.0577917
R848 VDD.n227 VDD.n226 0.0577917
R849 VDD.n237 VDD.n236 0.0577917
R850 VDD.n255 VDD.n254 0.0577917
R851 VDD.n265 VDD.n264 0.0577917
R852 VDD.n283 VDD.n282 0.0577917
R853 VDD.n293 VDD.n292 0.0577917
R854 VDD.n311 VDD.n310 0.0577917
R855 VDD.n321 VDD.n320 0.0577917
R856 VDD.n339 VDD.n338 0.0577917
R857 VDD.n349 VDD.n348 0.0577917
R858 VDD.n367 VDD.n366 0.0577917
R859 VDD.n377 VDD.n376 0.0577917
R860 VDD.n395 VDD.n394 0.0577917
R861 VDD.n405 VDD.n404 0.0577917
R862 VDD.n441 VDD.n422 0.0577917
R863 VDD.n436 VDD.n426 0.0577917
R864 VDD VDD.n211 0.00701042
R865 VDD VDD.n239 0.00701042
R866 VDD VDD.n267 0.00701042
R867 VDD VDD.n295 0.00701042
R868 VDD VDD.n323 0.00701042
R869 VDD VDD.n351 0.00701042
R870 VDD VDD.n379 0.00701042
R871 VDD.n456 VDD 0.00701042
R872 variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_unit_5.tristate_inverter_1.en.t7 628.097
R873 variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_unit_5.tristate_inverter_1.en.t2 622.766
R874 variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_unit_5.tristate_inverter_1.en.t5 523.774
R875 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t3 304.647
R876 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t4 304.647
R877 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t6 202.44
R878 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n0 168.969
R879 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n4 166.147
R880 variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_unit_5.tristate_inverter_1.en.t1 84.7557
R881 variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_unit_5.tristate_inverter_1.en.t0 84.1197
R882 variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_unit_5.tristate_inverter_1.en.n1 12.6535
R883 variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_unit_5.tristate_inverter_1.en 5.58443
R884 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n2 4.59003
R885 variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_unit_5.tristate_inverter_1.en.n3 1.09595
R886 variable_delay_unit_8.tristate_inverter_1.en.n3 variable_delay_unit_8.tristate_inverter_1.en.t3 628.097
R887 variable_delay_unit_8.tristate_inverter_1.en.n4 variable_delay_unit_8.tristate_inverter_1.en.t5 622.766
R888 variable_delay_unit_8.tristate_inverter_1.en.n3 variable_delay_unit_8.tristate_inverter_1.en.t7 523.774
R889 variable_delay_unit_8.tristate_inverter_1.en.n0 variable_delay_unit_8.tristate_inverter_1.en.t6 304.647
R890 variable_delay_unit_8.tristate_inverter_1.en.n0 variable_delay_unit_8.tristate_inverter_1.en.t2 304.647
R891 variable_delay_unit_8.tristate_inverter_1.en.n0 variable_delay_unit_8.tristate_inverter_1.en.t4 202.44
R892 variable_delay_unit_8.tristate_inverter_1.en variable_delay_unit_8.tristate_inverter_1.en.n0 168.969
R893 variable_delay_unit_8.tristate_inverter_1.en variable_delay_unit_8.tristate_inverter_1.en.n4 166.147
R894 variable_delay_unit_8.tristate_inverter_1.en.n1 variable_delay_unit_8.tristate_inverter_1.en.t1 84.7557
R895 variable_delay_unit_8.tristate_inverter_1.en.n1 variable_delay_unit_8.tristate_inverter_1.en.t0 84.1197
R896 variable_delay_unit_8.tristate_inverter_1.en.n2 variable_delay_unit_8.tristate_inverter_1.en.n1 12.6535
R897 variable_delay_unit_8.tristate_inverter_1.en.n2 variable_delay_unit_8.tristate_inverter_1.en 5.58443
R898 variable_delay_unit_8.tristate_inverter_1.en variable_delay_unit_8.tristate_inverter_1.en.n2 4.59003
R899 variable_delay_unit_8.tristate_inverter_1.en.n4 variable_delay_unit_8.tristate_inverter_1.en.n3 1.09595
R900 VSS.n135 VSS.n112 50016.6
R901 VSS.n483 VSS.n482 23663.9
R902 VSS.n386 VSS.n22 23663.9
R903 VSS.n385 VSS.n384 23663.9
R904 VSS.n300 VSS.n52 23663.9
R905 VSS.n299 VSS.n298 23663.9
R906 VSS.n214 VSS.n82 23663.9
R907 VSS.n213 VSS.n212 23663.9
R908 VSS.n491 VSS.n484 23663.9
R909 VSS.n492 VSS.n491 22860.5
R910 VSS.n149 VSS.n112 14239.4
R911 VSS.n213 VSS.n111 14239.4
R912 VSS.n235 VSS.n82 14239.4
R913 VSS.n299 VSS.n81 14239.4
R914 VSS.n321 VSS.n52 14239.4
R915 VSS.n385 VSS.n51 14239.4
R916 VSS.n407 VSS.n22 14239.4
R917 VSS.n483 VSS.n21 14239.4
R918 VSS.n491 VSS.n490 14239.4
R919 VSS.n212 VSS.n112 10823.2
R920 VSS.n214 VSS.n213 10823.2
R921 VSS.n298 VSS.n82 10823.2
R922 VSS.n300 VSS.n299 10823.2
R923 VSS.n384 VSS.n52 10823.2
R924 VSS.n386 VSS.n385 10823.2
R925 VSS.n482 VSS.n22 10823.2
R926 VSS.n484 VSS.n483 10823.2
R927 VSS.n484 VSS.n20 10102.8
R928 VSS.n212 VSS.n211 10102.8
R929 VSS.n218 VSS.n214 10102.8
R930 VSS.n298 VSS.n297 10102.8
R931 VSS.n304 VSS.n300 10102.8
R932 VSS.n384 VSS.n383 10102.8
R933 VSS.n390 VSS.n386 10102.8
R934 VSS.n482 VSS.n481 10102.8
R935 VSS.n146 VSS.n145 2045.07
R936 VSS.n198 VSS.n197 2045.07
R937 VSS.n232 VSS.n231 2045.07
R938 VSS.n284 VSS.n283 2045.07
R939 VSS.n318 VSS.n317 2045.07
R940 VSS.n370 VSS.n369 2045.07
R941 VSS.n404 VSS.n403 2045.07
R942 VSS.n468 VSS.n467 2045.07
R943 VSS.n515 VSS.n514 2045.07
R944 VSS.n516 VSS.n5 1626.7
R945 VSS.n18 VSS.n5 1626.7
R946 VSS.n471 VSS.n465 1626.7
R947 VSS.n471 VSS.n464 1626.7
R948 VSS.n433 VSS.n24 1626.7
R949 VSS.n479 VSS.n24 1626.7
R950 VSS.n410 VSS.n39 1626.7
R951 VSS.n410 VSS.n38 1626.7
R952 VSS.n402 VSS.n40 1626.7
R953 VSS.n388 VSS.n40 1626.7
R954 VSS.n373 VSS.n367 1626.7
R955 VSS.n373 VSS.n366 1626.7
R956 VSS.n347 VSS.n54 1626.7
R957 VSS.n381 VSS.n54 1626.7
R958 VSS.n324 VSS.n69 1626.7
R959 VSS.n324 VSS.n68 1626.7
R960 VSS.n316 VSS.n70 1626.7
R961 VSS.n302 VSS.n70 1626.7
R962 VSS.n287 VSS.n281 1626.7
R963 VSS.n287 VSS.n280 1626.7
R964 VSS.n261 VSS.n84 1626.7
R965 VSS.n295 VSS.n84 1626.7
R966 VSS.n238 VSS.n99 1626.7
R967 VSS.n238 VSS.n98 1626.7
R968 VSS.n230 VSS.n100 1626.7
R969 VSS.n216 VSS.n100 1626.7
R970 VSS.n201 VSS.n195 1626.7
R971 VSS.n201 VSS.n194 1626.7
R972 VSS.n175 VSS.n114 1626.7
R973 VSS.n209 VSS.n114 1626.7
R974 VSS.n152 VSS.n129 1626.7
R975 VSS.n152 VSS.n128 1626.7
R976 VSS.n144 VSS.n130 1626.7
R977 VSS.n136 VSS.n130 1626.7
R978 VSS.n486 VSS.n6 1626.7
R979 VSS.n513 VSS.n6 1626.7
R980 VSS.n219 VSS.n218 1460.78
R981 VSS.n297 VSS.n83 1460.78
R982 VSS.n305 VSS.n304 1460.78
R983 VSS.n383 VSS.n53 1460.78
R984 VSS.n391 VSS.n390 1460.78
R985 VSS.n481 VSS.n23 1460.78
R986 VSS.n446 VSS.n20 1460.78
R987 VSS.n211 VSS.n113 1460.78
R988 VSS.n211 VSS.n210 1437.75
R989 VSS.n218 VSS.n217 1437.75
R990 VSS.n297 VSS.n296 1437.75
R991 VSS.n304 VSS.n303 1437.75
R992 VSS.n383 VSS.n382 1437.75
R993 VSS.n390 VSS.n389 1437.75
R994 VSS.n481 VSS.n480 1437.75
R995 VSS.n20 VSS.n19 1437.75
R996 VSS.n185 VSS.n111 1138.52
R997 VSS.n235 VSS.n234 1138.52
R998 VSS.n271 VSS.n81 1138.52
R999 VSS.n321 VSS.n320 1138.52
R1000 VSS.n357 VSS.n51 1138.52
R1001 VSS.n407 VSS.n406 1138.52
R1002 VSS.n443 VSS.n21 1138.52
R1003 VSS.n149 VSS.n148 1138.52
R1004 VSS.n490 VSS.n489 1138.52
R1005 VSS.n150 VSS.n149 1115.49
R1006 VSS.n199 VSS.n111 1115.49
R1007 VSS.n236 VSS.n235 1115.49
R1008 VSS.n285 VSS.n81 1115.49
R1009 VSS.n322 VSS.n321 1115.49
R1010 VSS.n371 VSS.n51 1115.49
R1011 VSS.n408 VSS.n407 1115.49
R1012 VSS.n469 VSS.n21 1115.49
R1013 VSS.n490 VSS.n487 1115.49
R1014 VSS.n165 VSS.n119 1058.19
R1015 VSS.n165 VSS.n118 1058.19
R1016 VSS.n162 VSS.n120 1058.19
R1017 VSS.n147 VSS.n120 1058.19
R1018 VSS.n187 VSS.n182 1058.19
R1019 VSS.n184 VSS.n182 1058.19
R1020 VSS.n220 VSS.n109 1058.19
R1021 VSS.n220 VSS.n108 1058.19
R1022 VSS.n248 VSS.n90 1058.19
R1023 VSS.n233 VSS.n90 1058.19
R1024 VSS.n251 VSS.n89 1058.19
R1025 VSS.n251 VSS.n88 1058.19
R1026 VSS.n273 VSS.n268 1058.19
R1027 VSS.n270 VSS.n268 1058.19
R1028 VSS.n306 VSS.n79 1058.19
R1029 VSS.n306 VSS.n78 1058.19
R1030 VSS.n334 VSS.n60 1058.19
R1031 VSS.n319 VSS.n60 1058.19
R1032 VSS.n337 VSS.n59 1058.19
R1033 VSS.n337 VSS.n58 1058.19
R1034 VSS.n359 VSS.n354 1058.19
R1035 VSS.n356 VSS.n354 1058.19
R1036 VSS.n392 VSS.n49 1058.19
R1037 VSS.n392 VSS.n48 1058.19
R1038 VSS.n420 VSS.n30 1058.19
R1039 VSS.n405 VSS.n30 1058.19
R1040 VSS.n423 VSS.n29 1058.19
R1041 VSS.n423 VSS.n28 1058.19
R1042 VSS.n457 VSS.n440 1058.19
R1043 VSS.n442 VSS.n440 1058.19
R1044 VSS.n447 VSS.n444 1058.19
R1045 VSS.n454 VSS.n444 1058.19
R1046 VSS.n493 VSS.n15 1058.19
R1047 VSS.n500 VSS.n15 1058.19
R1048 VSS.n503 VSS.n13 1058.19
R1049 VSS.n488 VSS.n13 1058.19
R1050 VSS.t98 VSS.n185 943.788
R1051 VSS.n186 VSS.t98 943.788
R1052 VSS.t118 VSS.n110 943.788
R1053 VSS.t118 VSS.n219 943.788
R1054 VSS.n234 VSS.t27 943.788
R1055 VSS.n249 VSS.t27 943.788
R1056 VSS.t42 VSS.n250 943.788
R1057 VSS.t42 VSS.n83 943.788
R1058 VSS.t22 VSS.n271 943.788
R1059 VSS.n272 VSS.t22 943.788
R1060 VSS.t10 VSS.n80 943.788
R1061 VSS.t10 VSS.n305 943.788
R1062 VSS.n320 VSS.t47 943.788
R1063 VSS.n335 VSS.t47 943.788
R1064 VSS.t125 VSS.n336 943.788
R1065 VSS.t125 VSS.n53 943.788
R1066 VSS.t65 VSS.n357 943.788
R1067 VSS.n358 VSS.t65 943.788
R1068 VSS.t143 VSS.n50 943.788
R1069 VSS.t143 VSS.n391 943.788
R1070 VSS.n406 VSS.t112 943.788
R1071 VSS.n421 VSS.t112 943.788
R1072 VSS.t159 VSS.n422 943.788
R1073 VSS.t159 VSS.n23 943.788
R1074 VSS.t102 VSS.n443 943.788
R1075 VSS.n456 VSS.t102 943.788
R1076 VSS.n455 VSS.t63 943.788
R1077 VSS.n446 VSS.t63 943.788
R1078 VSS.n148 VSS.t96 943.788
R1079 VSS.n163 VSS.t96 943.788
R1080 VSS.t75 VSS.n164 943.788
R1081 VSS.t75 VSS.n113 943.788
R1082 VSS.n489 VSS.t161 943.788
R1083 VSS.n502 VSS.t161 943.788
R1084 VSS.n501 VSS.t32 943.788
R1085 VSS.n492 VSS.t32 943.788
R1086 VSS.n135 VSS.t4 892.394
R1087 VSS.n145 VSS.t55 892.394
R1088 VSS.t153 VSS.n146 892.394
R1089 VSS.t77 VSS.n150 892.394
R1090 VSS.n210 VSS.t108 892.394
R1091 VSS.n197 VSS.t56 892.394
R1092 VSS.t39 VSS.n198 892.394
R1093 VSS.t137 VSS.n199 892.394
R1094 VSS.n217 VSS.t87 892.394
R1095 VSS.n231 VSS.t105 892.394
R1096 VSS.t154 VSS.n232 892.394
R1097 VSS.t61 VSS.n236 892.394
R1098 VSS.n296 VSS.t91 892.394
R1099 VSS.n283 VSS.t53 892.394
R1100 VSS.t24 VSS.n284 892.394
R1101 VSS.t40 VSS.n285 892.394
R1102 VSS.n303 VSS.t81 892.394
R1103 VSS.n317 VSS.t14 892.394
R1104 VSS.t21 VSS.n318 892.394
R1105 VSS.t17 VSS.n322 892.394
R1106 VSS.n382 VSS.t85 892.394
R1107 VSS.n369 VSS.t104 892.394
R1108 VSS.t95 VSS.n370 892.394
R1109 VSS.t141 VSS.n371 892.394
R1110 VSS.n389 VSS.t49 892.394
R1111 VSS.n403 VSS.t155 892.394
R1112 VSS.t46 VSS.n404 892.394
R1113 VSS.t145 VSS.n408 892.394
R1114 VSS.n480 VSS.t131 892.394
R1115 VSS.n467 VSS.t120 892.394
R1116 VSS.t29 VSS.n468 892.394
R1117 VSS.t57 VSS.n469 892.394
R1118 VSS.n19 VSS.t37 892.394
R1119 VSS.n515 VSS.t156 892.394
R1120 VSS.n514 VSS.t34 892.394
R1121 VSS.n487 VSS.t30 892.394
R1122 VSS.n186 VSS.n110 702.96
R1123 VSS.n250 VSS.n249 702.96
R1124 VSS.n272 VSS.n80 702.96
R1125 VSS.n336 VSS.n335 702.96
R1126 VSS.n358 VSS.n50 702.96
R1127 VSS.n422 VSS.n421 702.96
R1128 VSS.n456 VSS.n455 702.96
R1129 VSS.n164 VSS.n163 702.96
R1130 VSS.n502 VSS.n501 702.96
R1131 VSS.n138 VSS.t163 607.409
R1132 VSS.t4 VSS.t2 545.352
R1133 VSS.t0 VSS.t55 545.352
R1134 VSS.t73 VSS.t153 545.352
R1135 VSS.t71 VSS.t77 545.352
R1136 VSS.t100 VSS.t108 545.352
R1137 VSS.t56 VSS.t133 545.352
R1138 VSS.t151 VSS.t39 545.352
R1139 VSS.t135 VSS.t137 545.352
R1140 VSS.t87 VSS.t147 545.352
R1141 VSS.t25 VSS.t105 545.352
R1142 VSS.t157 VSS.t154 545.352
R1143 VSS.t51 VSS.t61 545.352
R1144 VSS.t89 VSS.t91 545.352
R1145 VSS.t53 VSS.t93 545.352
R1146 VSS.t79 VSS.t24 545.352
R1147 VSS.t12 VSS.t40 545.352
R1148 VSS.t81 VSS.t110 545.352
R1149 VSS.t129 VSS.t14 545.352
R1150 VSS.t69 VSS.t21 545.352
R1151 VSS.t19 VSS.t17 545.352
R1152 VSS.t127 VSS.t85 545.352
R1153 VSS.t104 VSS.t83 545.352
R1154 VSS.t139 VSS.t95 545.352
R1155 VSS.t67 VSS.t141 545.352
R1156 VSS.t49 VSS.t59 545.352
R1157 VSS.t8 VSS.t155 545.352
R1158 VSS.t15 VSS.t46 545.352
R1159 VSS.t149 VSS.t145 545.352
R1160 VSS.t116 VSS.t131 545.352
R1161 VSS.t120 VSS.t121 545.352
R1162 VSS.t6 VSS.t29 545.352
R1163 VSS.t44 VSS.t57 545.352
R1164 VSS.t37 VSS.t35 545.352
R1165 VSS.t123 VSS.t156 545.352
R1166 VSS.t106 VSS.t34 545.352
R1167 VSS.t30 VSS.t114 545.352
R1168 VSS.n138 VSS.t54 321.423
R1169 VSS.t2 VSS.n134 272.676
R1170 VSS.n134 VSS.t0 272.676
R1171 VSS.n151 VSS.t73 272.676
R1172 VSS.n151 VSS.t71 272.676
R1173 VSS.n196 VSS.t100 272.676
R1174 VSS.t133 VSS.n196 272.676
R1175 VSS.n200 VSS.t151 272.676
R1176 VSS.n200 VSS.t135 272.676
R1177 VSS.t147 VSS.n215 272.676
R1178 VSS.n215 VSS.t25 272.676
R1179 VSS.n237 VSS.t157 272.676
R1180 VSS.n237 VSS.t51 272.676
R1181 VSS.n282 VSS.t89 272.676
R1182 VSS.t93 VSS.n282 272.676
R1183 VSS.n286 VSS.t79 272.676
R1184 VSS.n286 VSS.t12 272.676
R1185 VSS.t110 VSS.n301 272.676
R1186 VSS.n301 VSS.t129 272.676
R1187 VSS.n323 VSS.t69 272.676
R1188 VSS.n323 VSS.t19 272.676
R1189 VSS.n368 VSS.t127 272.676
R1190 VSS.t83 VSS.n368 272.676
R1191 VSS.n372 VSS.t139 272.676
R1192 VSS.n372 VSS.t67 272.676
R1193 VSS.t59 VSS.n387 272.676
R1194 VSS.n387 VSS.t8 272.676
R1195 VSS.n409 VSS.t15 272.676
R1196 VSS.n409 VSS.t149 272.676
R1197 VSS.n466 VSS.t116 272.676
R1198 VSS.t121 VSS.n466 272.676
R1199 VSS.n470 VSS.t6 272.676
R1200 VSS.n470 VSS.t44 272.676
R1201 VSS.t35 VSS.n17 272.676
R1202 VSS.n17 VSS.t123 272.676
R1203 VSS.n485 VSS.t106 272.676
R1204 VSS.t114 VSS.n485 272.676
R1205 VSS.n184 VSS.n180 195
R1206 VSS.n185 VSS.n184 195
R1207 VSS.n188 VSS.n187 195
R1208 VSS.n187 VSS.n186 195
R1209 VSS.n108 VSS.n107 195
R1210 VSS.n110 VSS.n108 195
R1211 VSS.n109 VSS.n105 195
R1212 VSS.n219 VSS.n109 195
R1213 VSS.n233 VSS.n92 195
R1214 VSS.n234 VSS.n233 195
R1215 VSS.n248 VSS.n247 195
R1216 VSS.n249 VSS.n248 195
R1217 VSS.n88 VSS.n87 195
R1218 VSS.n250 VSS.n88 195
R1219 VSS.n89 VSS.n85 195
R1220 VSS.n89 VSS.n83 195
R1221 VSS.n270 VSS.n266 195
R1222 VSS.n271 VSS.n270 195
R1223 VSS.n274 VSS.n273 195
R1224 VSS.n273 VSS.n272 195
R1225 VSS.n78 VSS.n77 195
R1226 VSS.n80 VSS.n78 195
R1227 VSS.n79 VSS.n75 195
R1228 VSS.n305 VSS.n79 195
R1229 VSS.n319 VSS.n62 195
R1230 VSS.n320 VSS.n319 195
R1231 VSS.n334 VSS.n333 195
R1232 VSS.n335 VSS.n334 195
R1233 VSS.n58 VSS.n57 195
R1234 VSS.n336 VSS.n58 195
R1235 VSS.n59 VSS.n55 195
R1236 VSS.n59 VSS.n53 195
R1237 VSS.n356 VSS.n352 195
R1238 VSS.n357 VSS.n356 195
R1239 VSS.n360 VSS.n359 195
R1240 VSS.n359 VSS.n358 195
R1241 VSS.n48 VSS.n47 195
R1242 VSS.n50 VSS.n48 195
R1243 VSS.n49 VSS.n45 195
R1244 VSS.n391 VSS.n49 195
R1245 VSS.n405 VSS.n32 195
R1246 VSS.n406 VSS.n405 195
R1247 VSS.n420 VSS.n419 195
R1248 VSS.n421 VSS.n420 195
R1249 VSS.n28 VSS.n27 195
R1250 VSS.n422 VSS.n28 195
R1251 VSS.n29 VSS.n25 195
R1252 VSS.n29 VSS.n23 195
R1253 VSS.n442 VSS.n438 195
R1254 VSS.n443 VSS.n442 195
R1255 VSS.n458 VSS.n457 195
R1256 VSS.n457 VSS.n456 195
R1257 VSS.n454 VSS.n453 195
R1258 VSS.n455 VSS.n454 195
R1259 VSS.n448 VSS.n447 195
R1260 VSS.n447 VSS.n446 195
R1261 VSS.n147 VSS.n122 195
R1262 VSS.n148 VSS.n147 195
R1263 VSS.n162 VSS.n161 195
R1264 VSS.n163 VSS.n162 195
R1265 VSS.n118 VSS.n117 195
R1266 VSS.n164 VSS.n118 195
R1267 VSS.n119 VSS.n115 195
R1268 VSS.n119 VSS.n113 195
R1269 VSS.n488 VSS.n11 195
R1270 VSS.n489 VSS.n488 195
R1271 VSS.n504 VSS.n503 195
R1272 VSS.n503 VSS.n502 195
R1273 VSS.n500 VSS.n499 195
R1274 VSS.n501 VSS.n500 195
R1275 VSS.n494 VSS.n493 195
R1276 VSS.n493 VSS.n492 195
R1277 VSS VSS.n138 161.595
R1278 VSS.n189 VSS.n182 146.25
R1279 VSS.t98 VSS.n182 146.25
R1280 VSS.n221 VSS.n220 146.25
R1281 VSS.n220 VSS.t118 146.25
R1282 VSS.n246 VSS.n90 146.25
R1283 VSS.n90 VSS.t27 146.25
R1284 VSS.n252 VSS.n251 146.25
R1285 VSS.n251 VSS.t42 146.25
R1286 VSS.n275 VSS.n268 146.25
R1287 VSS.t22 VSS.n268 146.25
R1288 VSS.n307 VSS.n306 146.25
R1289 VSS.n306 VSS.t10 146.25
R1290 VSS.n332 VSS.n60 146.25
R1291 VSS.n60 VSS.t47 146.25
R1292 VSS.n338 VSS.n337 146.25
R1293 VSS.n337 VSS.t125 146.25
R1294 VSS.n361 VSS.n354 146.25
R1295 VSS.t65 VSS.n354 146.25
R1296 VSS.n393 VSS.n392 146.25
R1297 VSS.n392 VSS.t143 146.25
R1298 VSS.n418 VSS.n30 146.25
R1299 VSS.n30 VSS.t112 146.25
R1300 VSS.n424 VSS.n423 146.25
R1301 VSS.n423 VSS.t159 146.25
R1302 VSS.n459 VSS.n440 146.25
R1303 VSS.t102 VSS.n440 146.25
R1304 VSS.n445 VSS.n444 146.25
R1305 VSS.n444 VSS.t63 146.25
R1306 VSS.n160 VSS.n120 146.25
R1307 VSS.n120 VSS.t96 146.25
R1308 VSS.n166 VSS.n165 146.25
R1309 VSS.n165 VSS.t75 146.25
R1310 VSS.n137 VSS.n136 146.25
R1311 VSS.n136 VSS.n135 146.25
R1312 VSS.n144 VSS.n143 146.25
R1313 VSS.n145 VSS.n144 146.25
R1314 VSS.n128 VSS.n127 146.25
R1315 VSS.n146 VSS.n128 146.25
R1316 VSS.n129 VSS.n123 146.25
R1317 VSS.n150 VSS.n129 146.25
R1318 VSS.n209 VSS.n208 146.25
R1319 VSS.n210 VSS.n209 146.25
R1320 VSS.n206 VSS.n175 146.25
R1321 VSS.n197 VSS.n175 146.25
R1322 VSS.n194 VSS.n176 146.25
R1323 VSS.n198 VSS.n194 146.25
R1324 VSS.n195 VSS.n193 146.25
R1325 VSS.n199 VSS.n195 146.25
R1326 VSS.n216 VSS.n104 146.25
R1327 VSS.n217 VSS.n216 146.25
R1328 VSS.n230 VSS.n229 146.25
R1329 VSS.n231 VSS.n230 146.25
R1330 VSS.n98 VSS.n97 146.25
R1331 VSS.n232 VSS.n98 146.25
R1332 VSS.n99 VSS.n93 146.25
R1333 VSS.n236 VSS.n99 146.25
R1334 VSS.n295 VSS.n294 146.25
R1335 VSS.n296 VSS.n295 146.25
R1336 VSS.n292 VSS.n261 146.25
R1337 VSS.n283 VSS.n261 146.25
R1338 VSS.n280 VSS.n262 146.25
R1339 VSS.n284 VSS.n280 146.25
R1340 VSS.n281 VSS.n279 146.25
R1341 VSS.n285 VSS.n281 146.25
R1342 VSS.n302 VSS.n74 146.25
R1343 VSS.n303 VSS.n302 146.25
R1344 VSS.n316 VSS.n315 146.25
R1345 VSS.n317 VSS.n316 146.25
R1346 VSS.n68 VSS.n67 146.25
R1347 VSS.n318 VSS.n68 146.25
R1348 VSS.n69 VSS.n63 146.25
R1349 VSS.n322 VSS.n69 146.25
R1350 VSS.n381 VSS.n380 146.25
R1351 VSS.n382 VSS.n381 146.25
R1352 VSS.n378 VSS.n347 146.25
R1353 VSS.n369 VSS.n347 146.25
R1354 VSS.n366 VSS.n348 146.25
R1355 VSS.n370 VSS.n366 146.25
R1356 VSS.n367 VSS.n365 146.25
R1357 VSS.n371 VSS.n367 146.25
R1358 VSS.n388 VSS.n44 146.25
R1359 VSS.n389 VSS.n388 146.25
R1360 VSS.n402 VSS.n401 146.25
R1361 VSS.n403 VSS.n402 146.25
R1362 VSS.n38 VSS.n37 146.25
R1363 VSS.n404 VSS.n38 146.25
R1364 VSS.n39 VSS.n33 146.25
R1365 VSS.n408 VSS.n39 146.25
R1366 VSS.n479 VSS.n478 146.25
R1367 VSS.n480 VSS.n479 146.25
R1368 VSS.n476 VSS.n433 146.25
R1369 VSS.n467 VSS.n433 146.25
R1370 VSS.n464 VSS.n434 146.25
R1371 VSS.n468 VSS.n464 146.25
R1372 VSS.n465 VSS.n463 146.25
R1373 VSS.n469 VSS.n465 146.25
R1374 VSS.n505 VSS.n13 146.25
R1375 VSS.t161 VSS.n13 146.25
R1376 VSS.n498 VSS.n15 146.25
R1377 VSS.n15 VSS.t32 146.25
R1378 VSS.n18 VSS.n4 146.25
R1379 VSS.n19 VSS.n18 146.25
R1380 VSS.n517 VSS.n516 146.25
R1381 VSS.n516 VSS.n515 146.25
R1382 VSS.n513 VSS.n512 146.25
R1383 VSS.n514 VSS.n513 146.25
R1384 VSS.n486 VSS.n10 146.25
R1385 VSS.n487 VSS.n486 146.25
R1386 VSS.n518 VSS.n517 105.695
R1387 VSS.n518 VSS.n4 105.695
R1388 VSS.n208 VSS.n207 105.695
R1389 VSS.n207 VSS.n206 105.695
R1390 VSS.n202 VSS.n176 105.695
R1391 VSS.n202 VSS.n193 105.695
R1392 VSS.n104 VSS.n101 105.695
R1393 VSS.n229 VSS.n101 105.695
R1394 VSS.n239 VSS.n97 105.695
R1395 VSS.n239 VSS.n93 105.695
R1396 VSS.n294 VSS.n293 105.695
R1397 VSS.n293 VSS.n292 105.695
R1398 VSS.n288 VSS.n262 105.695
R1399 VSS.n288 VSS.n279 105.695
R1400 VSS.n74 VSS.n71 105.695
R1401 VSS.n315 VSS.n71 105.695
R1402 VSS.n325 VSS.n67 105.695
R1403 VSS.n325 VSS.n63 105.695
R1404 VSS.n380 VSS.n379 105.695
R1405 VSS.n379 VSS.n378 105.695
R1406 VSS.n374 VSS.n348 105.695
R1407 VSS.n374 VSS.n365 105.695
R1408 VSS.n44 VSS.n41 105.695
R1409 VSS.n401 VSS.n41 105.695
R1410 VSS.n411 VSS.n37 105.695
R1411 VSS.n411 VSS.n33 105.695
R1412 VSS.n478 VSS.n477 105.695
R1413 VSS.n477 VSS.n476 105.695
R1414 VSS.n472 VSS.n434 105.695
R1415 VSS.n472 VSS.n463 105.695
R1416 VSS.n137 VSS.n131 105.695
R1417 VSS.n143 VSS.n131 105.695
R1418 VSS.n153 VSS.n127 105.695
R1419 VSS.n153 VSS.n123 105.695
R1420 VSS.n512 VSS.n7 105.695
R1421 VSS.n10 VSS.n7 105.695
R1422 VSS.n12 VSS.t162 84.1574
R1423 VSS.n496 VSS.t33 84.1574
R1424 VSS.n158 VSS.t97 84.1574
R1425 VSS.n168 VSS.t76 84.1574
R1426 VSS.n181 VSS.t99 84.1574
R1427 VSS.n223 VSS.t119 84.1574
R1428 VSS.n244 VSS.t28 84.1574
R1429 VSS.n254 VSS.t43 84.1574
R1430 VSS.n267 VSS.t23 84.1574
R1431 VSS.n309 VSS.t11 84.1574
R1432 VSS.n330 VSS.t48 84.1574
R1433 VSS.n340 VSS.t126 84.1574
R1434 VSS.n353 VSS.t66 84.1574
R1435 VSS.n395 VSS.t144 84.1574
R1436 VSS.n416 VSS.t113 84.1574
R1437 VSS.n426 VSS.t160 84.1574
R1438 VSS.n439 VSS.t103 84.1574
R1439 VSS.n450 VSS.t64 84.1574
R1440 VSS.n2 VSS.t38 83.7172
R1441 VSS.n9 VSS.t31 83.7172
R1442 VSS.n172 VSS.t109 83.7172
R1443 VSS.n178 VSS.t138 83.7172
R1444 VSS.n103 VSS.t88 83.7172
R1445 VSS.n95 VSS.t62 83.7172
R1446 VSS.n258 VSS.t92 83.7172
R1447 VSS.n264 VSS.t41 83.7172
R1448 VSS.n73 VSS.t82 83.7172
R1449 VSS.n65 VSS.t18 83.7172
R1450 VSS.n344 VSS.t86 83.7172
R1451 VSS.n350 VSS.t142 83.7172
R1452 VSS.n43 VSS.t50 83.7172
R1453 VSS.n35 VSS.t146 83.7172
R1454 VSS.n430 VSS.t132 83.7172
R1455 VSS.n436 VSS.t58 83.7172
R1456 VSS.n133 VSS.t5 83.7172
R1457 VSS.n125 VSS.t78 83.7172
R1458 VSS.n2 VSS.n1 75.905
R1459 VSS.n9 VSS.n8 75.905
R1460 VSS.n172 VSS.n171 75.905
R1461 VSS.n178 VSS.n177 75.905
R1462 VSS.n103 VSS.n102 75.905
R1463 VSS.n95 VSS.n94 75.905
R1464 VSS.n258 VSS.n257 75.905
R1465 VSS.n264 VSS.n263 75.905
R1466 VSS.n73 VSS.n72 75.905
R1467 VSS.n65 VSS.n64 75.905
R1468 VSS.n344 VSS.n343 75.905
R1469 VSS.n350 VSS.n349 75.905
R1470 VSS.n43 VSS.n42 75.905
R1471 VSS.n35 VSS.n34 75.905
R1472 VSS.n430 VSS.n429 75.905
R1473 VSS.n436 VSS.n435 75.905
R1474 VSS.n133 VSS.n132 75.905
R1475 VSS.n125 VSS.n124 75.905
R1476 VSS.n131 VSS.n130 73.1255
R1477 VSS.n134 VSS.n130 73.1255
R1478 VSS.n153 VSS.n152 73.1255
R1479 VSS.n152 VSS.n151 73.1255
R1480 VSS.n207 VSS.n114 73.1255
R1481 VSS.n196 VSS.n114 73.1255
R1482 VSS.n202 VSS.n201 73.1255
R1483 VSS.n201 VSS.n200 73.1255
R1484 VSS.n101 VSS.n100 73.1255
R1485 VSS.n215 VSS.n100 73.1255
R1486 VSS.n239 VSS.n238 73.1255
R1487 VSS.n238 VSS.n237 73.1255
R1488 VSS.n293 VSS.n84 73.1255
R1489 VSS.n282 VSS.n84 73.1255
R1490 VSS.n288 VSS.n287 73.1255
R1491 VSS.n287 VSS.n286 73.1255
R1492 VSS.n71 VSS.n70 73.1255
R1493 VSS.n301 VSS.n70 73.1255
R1494 VSS.n325 VSS.n324 73.1255
R1495 VSS.n324 VSS.n323 73.1255
R1496 VSS.n379 VSS.n54 73.1255
R1497 VSS.n368 VSS.n54 73.1255
R1498 VSS.n374 VSS.n373 73.1255
R1499 VSS.n373 VSS.n372 73.1255
R1500 VSS.n41 VSS.n40 73.1255
R1501 VSS.n387 VSS.n40 73.1255
R1502 VSS.n411 VSS.n410 73.1255
R1503 VSS.n410 VSS.n409 73.1255
R1504 VSS.n477 VSS.n24 73.1255
R1505 VSS.n466 VSS.n24 73.1255
R1506 VSS.n472 VSS.n471 73.1255
R1507 VSS.n471 VSS.n470 73.1255
R1508 VSS.n518 VSS.n5 73.1255
R1509 VSS.n17 VSS.n5 73.1255
R1510 VSS.n7 VSS.n6 73.1255
R1511 VSS.n485 VSS.n6 73.1255
R1512 VSS.n166 VSS.n117 68.7561
R1513 VSS.n166 VSS.n115 68.7561
R1514 VSS.n189 VSS.n188 68.7561
R1515 VSS.n189 VSS.n180 68.7561
R1516 VSS.n221 VSS.n107 68.7561
R1517 VSS.n221 VSS.n105 68.7561
R1518 VSS.n247 VSS.n246 68.7561
R1519 VSS.n246 VSS.n92 68.7561
R1520 VSS.n252 VSS.n87 68.7561
R1521 VSS.n252 VSS.n85 68.7561
R1522 VSS.n275 VSS.n274 68.7561
R1523 VSS.n275 VSS.n266 68.7561
R1524 VSS.n307 VSS.n77 68.7561
R1525 VSS.n307 VSS.n75 68.7561
R1526 VSS.n333 VSS.n332 68.7561
R1527 VSS.n332 VSS.n62 68.7561
R1528 VSS.n338 VSS.n57 68.7561
R1529 VSS.n338 VSS.n55 68.7561
R1530 VSS.n361 VSS.n360 68.7561
R1531 VSS.n361 VSS.n352 68.7561
R1532 VSS.n393 VSS.n47 68.7561
R1533 VSS.n393 VSS.n45 68.7561
R1534 VSS.n419 VSS.n418 68.7561
R1535 VSS.n418 VSS.n32 68.7561
R1536 VSS.n424 VSS.n27 68.7561
R1537 VSS.n424 VSS.n25 68.7561
R1538 VSS.n459 VSS.n458 68.7561
R1539 VSS.n459 VSS.n438 68.7561
R1540 VSS.n453 VSS.n445 68.7561
R1541 VSS.n448 VSS.n445 68.7561
R1542 VSS.n161 VSS.n160 68.7561
R1543 VSS.n160 VSS.n122 68.7561
R1544 VSS.n498 VSS.n494 68.7561
R1545 VSS.n499 VSS.n498 68.7561
R1546 VSS.n505 VSS.n504 68.7561
R1547 VSS.n505 VSS.n11 68.7561
R1548 VSS.n1 VSS.t36 17.4005
R1549 VSS.n1 VSS.t124 17.4005
R1550 VSS.n8 VSS.t107 17.4005
R1551 VSS.n8 VSS.t115 17.4005
R1552 VSS.n171 VSS.t101 17.4005
R1553 VSS.n171 VSS.t134 17.4005
R1554 VSS.n177 VSS.t152 17.4005
R1555 VSS.n177 VSS.t136 17.4005
R1556 VSS.n102 VSS.t148 17.4005
R1557 VSS.n102 VSS.t26 17.4005
R1558 VSS.n94 VSS.t158 17.4005
R1559 VSS.n94 VSS.t52 17.4005
R1560 VSS.n257 VSS.t90 17.4005
R1561 VSS.n257 VSS.t94 17.4005
R1562 VSS.n263 VSS.t80 17.4005
R1563 VSS.n263 VSS.t13 17.4005
R1564 VSS.n72 VSS.t111 17.4005
R1565 VSS.n72 VSS.t130 17.4005
R1566 VSS.n64 VSS.t70 17.4005
R1567 VSS.n64 VSS.t20 17.4005
R1568 VSS.n343 VSS.t128 17.4005
R1569 VSS.n343 VSS.t84 17.4005
R1570 VSS.n349 VSS.t140 17.4005
R1571 VSS.n349 VSS.t68 17.4005
R1572 VSS.n42 VSS.t60 17.4005
R1573 VSS.n42 VSS.t9 17.4005
R1574 VSS.n34 VSS.t16 17.4005
R1575 VSS.n34 VSS.t150 17.4005
R1576 VSS.n429 VSS.t117 17.4005
R1577 VSS.n429 VSS.t122 17.4005
R1578 VSS.n435 VSS.t7 17.4005
R1579 VSS.n435 VSS.t45 17.4005
R1580 VSS.n132 VSS.t3 17.4005
R1581 VSS.n132 VSS.t1 17.4005
R1582 VSS.n124 VSS.t74 17.4005
R1583 VSS.n124 VSS.t72 17.4005
R1584 VSS.n157 VSS.n122 3.46248
R1585 VSS.n117 VSS.n116 3.46248
R1586 VSS.n169 VSS.n115 3.46248
R1587 VSS.n107 VSS.n106 3.46248
R1588 VSS.n191 VSS.n180 3.46248
R1589 VSS.n188 VSS.n183 3.46248
R1590 VSS.n224 VSS.n105 3.46248
R1591 VSS.n87 VSS.n86 3.46248
R1592 VSS.n243 VSS.n92 3.46248
R1593 VSS.n247 VSS.n91 3.46248
R1594 VSS.n255 VSS.n85 3.46248
R1595 VSS.n77 VSS.n76 3.46248
R1596 VSS.n277 VSS.n266 3.46248
R1597 VSS.n274 VSS.n269 3.46248
R1598 VSS.n310 VSS.n75 3.46248
R1599 VSS.n57 VSS.n56 3.46248
R1600 VSS.n329 VSS.n62 3.46248
R1601 VSS.n333 VSS.n61 3.46248
R1602 VSS.n341 VSS.n55 3.46248
R1603 VSS.n47 VSS.n46 3.46248
R1604 VSS.n363 VSS.n352 3.46248
R1605 VSS.n360 VSS.n355 3.46248
R1606 VSS.n396 VSS.n45 3.46248
R1607 VSS.n27 VSS.n26 3.46248
R1608 VSS.n415 VSS.n32 3.46248
R1609 VSS.n419 VSS.n31 3.46248
R1610 VSS.n427 VSS.n25 3.46248
R1611 VSS.n453 VSS.n452 3.46248
R1612 VSS.n461 VSS.n438 3.46248
R1613 VSS.n458 VSS.n441 3.46248
R1614 VSS.n449 VSS.n448 3.46248
R1615 VSS.n161 VSS.n121 3.46248
R1616 VSS.n499 VSS.n16 3.46248
R1617 VSS.n495 VSS.n494 3.46248
R1618 VSS.n507 VSS.n11 3.46248
R1619 VSS.n504 VSS.n14 3.46248
R1620 VSS.n512 VSS.n511 2.82278
R1621 VSS.n4 VSS.n0 2.82278
R1622 VSS.n517 VSS.n3 2.82278
R1623 VSS.n208 VSS.n170 2.82278
R1624 VSS.n206 VSS.n205 2.82278
R1625 VSS.n204 VSS.n176 2.82278
R1626 VSS.n193 VSS.n192 2.82278
R1627 VSS.n225 VSS.n104 2.82278
R1628 VSS.n229 VSS.n228 2.82278
R1629 VSS.n97 VSS.n96 2.82278
R1630 VSS.n242 VSS.n93 2.82278
R1631 VSS.n294 VSS.n256 2.82278
R1632 VSS.n292 VSS.n291 2.82278
R1633 VSS.n290 VSS.n262 2.82278
R1634 VSS.n279 VSS.n278 2.82278
R1635 VSS.n311 VSS.n74 2.82278
R1636 VSS.n315 VSS.n314 2.82278
R1637 VSS.n67 VSS.n66 2.82278
R1638 VSS.n328 VSS.n63 2.82278
R1639 VSS.n380 VSS.n342 2.82278
R1640 VSS.n378 VSS.n377 2.82278
R1641 VSS.n376 VSS.n348 2.82278
R1642 VSS.n365 VSS.n364 2.82278
R1643 VSS.n397 VSS.n44 2.82278
R1644 VSS.n401 VSS.n400 2.82278
R1645 VSS.n37 VSS.n36 2.82278
R1646 VSS.n414 VSS.n33 2.82278
R1647 VSS.n478 VSS.n428 2.82278
R1648 VSS.n476 VSS.n475 2.82278
R1649 VSS.n474 VSS.n434 2.82278
R1650 VSS.n463 VSS.n462 2.82278
R1651 VSS.n139 VSS.n137 2.82278
R1652 VSS.n143 VSS.n142 2.82278
R1653 VSS.n127 VSS.n126 2.82278
R1654 VSS.n156 VSS.n123 2.82278
R1655 VSS.n508 VSS.n10 2.82278
R1656 VSS.n460 VSS.n459 2.3255
R1657 VSS.n451 VSS.n445 2.3255
R1658 VSS.n418 VSS.n417 2.3255
R1659 VSS.n425 VSS.n424 2.3255
R1660 VSS.n362 VSS.n361 2.3255
R1661 VSS.n394 VSS.n393 2.3255
R1662 VSS.n332 VSS.n331 2.3255
R1663 VSS.n339 VSS.n338 2.3255
R1664 VSS.n276 VSS.n275 2.3255
R1665 VSS.n308 VSS.n307 2.3255
R1666 VSS.n246 VSS.n245 2.3255
R1667 VSS.n253 VSS.n252 2.3255
R1668 VSS.n190 VSS.n189 2.3255
R1669 VSS.n222 VSS.n221 2.3255
R1670 VSS.n167 VSS.n166 2.3255
R1671 VSS.n160 VSS.n159 2.3255
R1672 VSS.n506 VSS.n505 2.3255
R1673 VSS.n498 VSS.n497 2.3255
R1674 VSS.n477 VSS.n432 1.32907
R1675 VSS.n473 VSS.n472 1.32907
R1676 VSS.n399 VSS.n41 1.32907
R1677 VSS.n412 VSS.n411 1.32907
R1678 VSS.n379 VSS.n346 1.32907
R1679 VSS.n375 VSS.n374 1.32907
R1680 VSS.n313 VSS.n71 1.32907
R1681 VSS.n326 VSS.n325 1.32907
R1682 VSS.n293 VSS.n260 1.32907
R1683 VSS.n289 VSS.n288 1.32907
R1684 VSS.n227 VSS.n101 1.32907
R1685 VSS.n240 VSS.n239 1.32907
R1686 VSS.n207 VSS.n174 1.32907
R1687 VSS.n203 VSS.n202 1.32907
R1688 VSS.n141 VSS.n131 1.32907
R1689 VSS.n154 VSS.n153 1.32907
R1690 VSS.n519 VSS.n518 1.32907
R1691 VSS.n510 VSS.n7 1.32907
R1692 VSS.n139 VSS 1.14229
R1693 VSS.n520 VSS.n2 0.685283
R1694 VSS.n509 VSS.n9 0.685283
R1695 VSS.n173 VSS.n172 0.685283
R1696 VSS.n179 VSS.n178 0.685283
R1697 VSS.n226 VSS.n103 0.685283
R1698 VSS.n241 VSS.n95 0.685283
R1699 VSS.n259 VSS.n258 0.685283
R1700 VSS.n265 VSS.n264 0.685283
R1701 VSS.n312 VSS.n73 0.685283
R1702 VSS.n327 VSS.n65 0.685283
R1703 VSS.n345 VSS.n344 0.685283
R1704 VSS.n351 VSS.n350 0.685283
R1705 VSS.n398 VSS.n43 0.685283
R1706 VSS.n413 VSS.n35 0.685283
R1707 VSS.n431 VSS.n430 0.685283
R1708 VSS.n437 VSS.n436 0.685283
R1709 VSS.n140 VSS.n133 0.685283
R1710 VSS.n155 VSS.n125 0.685283
R1711 VSS.n449 VSS 0.479667
R1712 VSS VSS.n427 0.479667
R1713 VSS VSS.n396 0.479667
R1714 VSS VSS.n341 0.479667
R1715 VSS VSS.n310 0.479667
R1716 VSS VSS.n255 0.479667
R1717 VSS VSS.n224 0.479667
R1718 VSS VSS.n169 0.479667
R1719 VSS VSS.n461 0.466646
R1720 VSS.n415 VSS 0.466646
R1721 VSS VSS.n363 0.466646
R1722 VSS.n329 VSS 0.466646
R1723 VSS VSS.n277 0.466646
R1724 VSS.n243 VSS 0.466646
R1725 VSS VSS.n191 0.466646
R1726 VSS.n157 VSS 0.466646
R1727 VSS VSS.n507 0.466646
R1728 VSS.n475 VSS.n474 0.430188
R1729 VSS.n400 VSS.n36 0.430188
R1730 VSS.n377 VSS.n376 0.430188
R1731 VSS.n314 VSS.n66 0.430188
R1732 VSS.n291 VSS.n290 0.430188
R1733 VSS.n228 VSS.n96 0.430188
R1734 VSS.n205 VSS.n204 0.430188
R1735 VSS.n142 VSS.n126 0.430188
R1736 VSS.n511 VSS.n3 0.430188
R1737 VSS.n495 VSS 0.404146
R1738 VSS.n475 VSS.n432 0.359875
R1739 VSS.n474 VSS.n473 0.359875
R1740 VSS.n400 VSS.n399 0.359875
R1741 VSS.n412 VSS.n36 0.359875
R1742 VSS.n377 VSS.n346 0.359875
R1743 VSS.n376 VSS.n375 0.359875
R1744 VSS.n314 VSS.n313 0.359875
R1745 VSS.n326 VSS.n66 0.359875
R1746 VSS.n291 VSS.n260 0.359875
R1747 VSS.n290 VSS.n289 0.359875
R1748 VSS.n228 VSS.n227 0.359875
R1749 VSS.n240 VSS.n96 0.359875
R1750 VSS.n205 VSS.n174 0.359875
R1751 VSS.n204 VSS.n203 0.359875
R1752 VSS.n142 VSS.n141 0.359875
R1753 VSS.n154 VSS.n126 0.359875
R1754 VSS.n519 VSS.n3 0.359875
R1755 VSS.n511 VSS.n510 0.359875
R1756 VSS.n432 VSS.n431 0.229667
R1757 VSS.n473 VSS.n437 0.229667
R1758 VSS.n399 VSS.n398 0.229667
R1759 VSS.n413 VSS.n412 0.229667
R1760 VSS.n346 VSS.n345 0.229667
R1761 VSS.n375 VSS.n351 0.229667
R1762 VSS.n313 VSS.n312 0.229667
R1763 VSS.n327 VSS.n326 0.229667
R1764 VSS.n260 VSS.n259 0.229667
R1765 VSS.n289 VSS.n265 0.229667
R1766 VSS.n227 VSS.n226 0.229667
R1767 VSS.n241 VSS.n240 0.229667
R1768 VSS.n174 VSS.n173 0.229667
R1769 VSS.n203 VSS.n179 0.229667
R1770 VSS.n141 VSS.n140 0.229667
R1771 VSS.n155 VSS.n154 0.229667
R1772 VSS.n520 VSS.n519 0.229667
R1773 VSS.n510 VSS.n509 0.229667
R1774 VSS.n428 VSS 0.191906
R1775 VSS.n397 VSS 0.191906
R1776 VSS.n342 VSS 0.191906
R1777 VSS.n311 VSS 0.191906
R1778 VSS.n256 VSS 0.191906
R1779 VSS.n225 VSS 0.191906
R1780 VSS.n170 VSS 0.191906
R1781 VSS VSS.n0 0.191906
R1782 VSS.n461 VSS.n460 0.189302
R1783 VSS.n452 VSS.n451 0.189302
R1784 VSS.n417 VSS.n415 0.189302
R1785 VSS.n425 VSS.n26 0.189302
R1786 VSS.n363 VSS.n362 0.189302
R1787 VSS.n394 VSS.n46 0.189302
R1788 VSS.n331 VSS.n329 0.189302
R1789 VSS.n339 VSS.n56 0.189302
R1790 VSS.n277 VSS.n276 0.189302
R1791 VSS.n308 VSS.n76 0.189302
R1792 VSS.n245 VSS.n243 0.189302
R1793 VSS.n253 VSS.n86 0.189302
R1794 VSS.n191 VSS.n190 0.189302
R1795 VSS.n222 VSS.n106 0.189302
R1796 VSS.n159 VSS.n157 0.189302
R1797 VSS.n167 VSS.n116 0.189302
R1798 VSS.n507 VSS.n506 0.189302
R1799 VSS.n497 VSS.n16 0.189302
R1800 VSS.n452 VSS.n441 0.141125
R1801 VSS.n31 VSS.n26 0.141125
R1802 VSS.n355 VSS.n46 0.141125
R1803 VSS.n61 VSS.n56 0.141125
R1804 VSS.n269 VSS.n76 0.141125
R1805 VSS.n91 VSS.n86 0.141125
R1806 VSS.n183 VSS.n106 0.141125
R1807 VSS.n121 VSS.n116 0.141125
R1808 VSS.n16 VSS.n14 0.141125
R1809 VSS.n441 VSS.n439 0.13201
R1810 VSS.n450 VSS.n449 0.13201
R1811 VSS.n416 VSS.n31 0.13201
R1812 VSS.n427 VSS.n426 0.13201
R1813 VSS.n355 VSS.n353 0.13201
R1814 VSS.n396 VSS.n395 0.13201
R1815 VSS.n330 VSS.n61 0.13201
R1816 VSS.n341 VSS.n340 0.13201
R1817 VSS.n269 VSS.n267 0.13201
R1818 VSS.n310 VSS.n309 0.13201
R1819 VSS.n244 VSS.n91 0.13201
R1820 VSS.n255 VSS.n254 0.13201
R1821 VSS.n183 VSS.n181 0.13201
R1822 VSS.n224 VSS.n223 0.13201
R1823 VSS.n158 VSS.n121 0.13201
R1824 VSS.n169 VSS.n168 0.13201
R1825 VSS.n14 VSS.n12 0.13201
R1826 VSS.n496 VSS.n495 0.13201
R1827 VSS.n462 VSS.n437 0.130708
R1828 VSS.n414 VSS.n413 0.130708
R1829 VSS.n364 VSS.n351 0.130708
R1830 VSS.n328 VSS.n327 0.130708
R1831 VSS.n278 VSS.n265 0.130708
R1832 VSS.n242 VSS.n241 0.130708
R1833 VSS.n192 VSS.n179 0.130708
R1834 VSS.n156 VSS.n155 0.130708
R1835 VSS.n509 VSS.n508 0.130708
R1836 VSS.n431 VSS 0.124198
R1837 VSS.n398 VSS 0.124198
R1838 VSS.n345 VSS 0.124198
R1839 VSS.n312 VSS 0.124198
R1840 VSS.n259 VSS 0.124198
R1841 VSS.n226 VSS 0.124198
R1842 VSS.n173 VSS 0.124198
R1843 VSS.n140 VSS 0.124198
R1844 VSS VSS.n520 0.124198
R1845 VSS.n462 VSS 0.0695104
R1846 VSS VSS.n414 0.0695104
R1847 VSS.n364 VSS 0.0695104
R1848 VSS VSS.n328 0.0695104
R1849 VSS.n278 VSS 0.0695104
R1850 VSS VSS.n242 0.0695104
R1851 VSS.n192 VSS 0.0695104
R1852 VSS VSS.n156 0.0695104
R1853 VSS.n508 VSS 0.0695104
R1854 VSS.n460 VSS.n439 0.0577917
R1855 VSS.n451 VSS.n450 0.0577917
R1856 VSS.n417 VSS.n416 0.0577917
R1857 VSS.n426 VSS.n425 0.0577917
R1858 VSS.n362 VSS.n353 0.0577917
R1859 VSS.n395 VSS.n394 0.0577917
R1860 VSS.n331 VSS.n330 0.0577917
R1861 VSS.n340 VSS.n339 0.0577917
R1862 VSS.n276 VSS.n267 0.0577917
R1863 VSS.n309 VSS.n308 0.0577917
R1864 VSS.n245 VSS.n244 0.0577917
R1865 VSS.n254 VSS.n253 0.0577917
R1866 VSS.n190 VSS.n181 0.0577917
R1867 VSS.n223 VSS.n222 0.0577917
R1868 VSS.n159 VSS.n158 0.0577917
R1869 VSS.n168 VSS.n167 0.0577917
R1870 VSS.n506 VSS.n12 0.0577917
R1871 VSS.n497 VSS.n496 0.0577917
R1872 VSS VSS.n428 0.00701042
R1873 VSS VSS.n397 0.00701042
R1874 VSS VSS.n342 0.00701042
R1875 VSS VSS.n311 0.00701042
R1876 VSS VSS.n256 0.00701042
R1877 VSS VSS.n225 0.00701042
R1878 VSS VSS.n170 0.00701042
R1879 VSS VSS.n139 0.00701042
R1880 VSS VSS.n0 0.00701042
R1881 en_6.n0 en_6.t5 628.097
R1882 en_6.n1 en_6.t3 622.766
R1883 en_6.n2 en_6.t6 543.053
R1884 en_6.n0 en_6.t1 523.774
R1885 en_6.n4 en_6.t4 304.647
R1886 en_6.n4 en_6.t0 304.647
R1887 en_6.n2 en_6.t7 221.72
R1888 en_6 en_6.n2 220.304
R1889 en_6.n4 en_6.t2 202.44
R1890 en_6 en_6.n4 168.969
R1891 en_6 en_6.n1 166.147
R1892 en_6.n3 en_6 3.22371
R1893 en_6.n3 en_6 1.40175
R1894 en_6.n1 en_6.n0 1.09595
R1895 en_6 en_6.n3 0.443357
R1896 en_1.n2 en_1.t0 628.097
R1897 en_1.n3 en_1.t1 622.766
R1898 en_1.n0 en_1.t4 543.053
R1899 en_1.n2 en_1.t3 523.774
R1900 en_1.n1 en_1.t6 304.647
R1901 en_1.n1 en_1.t7 304.647
R1902 en_1.n0 en_1.t5 221.72
R1903 en_1.n5 en_1.n0 220.263
R1904 en_1.n1 en_1.t2 202.44
R1905 en_1 en_1.n1 168.969
R1906 en_1 en_1.n3 166.147
R1907 en_1 en_1.n4 3.15943
R1908 en_1.n4 en_1 1.40175
R1909 en_1.n3 en_1.n2 1.09595
R1910 en_1.n4 en_1 0.443357
R1911 en_1.n5 en_1 0.105857
R1912 en_1 en_1.n5 0.063
R1913 variable_delay_unit_3.in.n0 variable_delay_unit_3.in.t4 607.409
R1914 variable_delay_unit_3.in.n2 variable_delay_unit_3.in.t2 543.053
R1915 variable_delay_unit_3.in.n0 variable_delay_unit_3.in.t5 321.423
R1916 variable_delay_unit_3.in variable_delay_unit_3.in.n2 221.778
R1917 variable_delay_unit_3.in.n2 variable_delay_unit_3.in.t3 221.72
R1918 variable_delay_unit_3.in variable_delay_unit_3.in.n0 161.72
R1919 variable_delay_unit_3.in.n1 variable_delay_unit_3.in.t0 84.7227
R1920 variable_delay_unit_3.in.n1 variable_delay_unit_3.in.t1 84.0867
R1921 variable_delay_unit_3.in.n3 variable_delay_unit_3.in 20.0791
R1922 variable_delay_unit_3.in variable_delay_unit_3.in.n3 0.851271
R1923 variable_delay_unit_3.in.n3 variable_delay_unit_3.in.n1 0.465495
R1924 variable_delay_unit_4.in.n0 variable_delay_unit_4.in.t3 607.409
R1925 variable_delay_unit_4.in.n2 variable_delay_unit_4.in.t2 543.053
R1926 variable_delay_unit_4.in.n0 variable_delay_unit_4.in.t5 321.423
R1927 variable_delay_unit_4.in variable_delay_unit_4.in.n2 221.778
R1928 variable_delay_unit_4.in.n2 variable_delay_unit_4.in.t4 221.72
R1929 variable_delay_unit_4.in variable_delay_unit_4.in.n0 161.72
R1930 variable_delay_unit_4.in.n1 variable_delay_unit_4.in.t1 84.7227
R1931 variable_delay_unit_4.in.n1 variable_delay_unit_4.in.t0 84.0867
R1932 variable_delay_unit_4.in.n3 variable_delay_unit_4.in 20.0791
R1933 variable_delay_unit_4.in variable_delay_unit_4.in.n3 0.851271
R1934 variable_delay_unit_4.in.n3 variable_delay_unit_4.in.n1 0.465495
R1935 variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_unit_2.tristate_inverter_1.en.t5 628.097
R1936 variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_unit_2.tristate_inverter_1.en.t7 622.766
R1937 variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_unit_2.tristate_inverter_1.en.t3 523.774
R1938 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t2 304.647
R1939 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t4 304.647
R1940 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t6 202.44
R1941 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n0 168.969
R1942 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n4 166.147
R1943 variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_unit_2.tristate_inverter_1.en.t1 84.7557
R1944 variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_unit_2.tristate_inverter_1.en.t0 84.1197
R1945 variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_unit_2.tristate_inverter_1.en.n1 12.6535
R1946 variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_unit_2.tristate_inverter_1.en 5.58443
R1947 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n2 4.59003
R1948 variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_unit_2.tristate_inverter_1.en.n3 1.09595
R1949 variable_delay_unit_8.forward.n0 variable_delay_unit_8.forward.t2 607.409
R1950 variable_delay_unit_8.forward.n0 variable_delay_unit_8.forward.t3 321.423
R1951 variable_delay_unit_8.forward variable_delay_unit_8.forward.n0 161.72
R1952 variable_delay_unit_8.forward.n1 variable_delay_unit_8.forward.t1 84.7227
R1953 variable_delay_unit_8.forward.n1 variable_delay_unit_8.forward.t0 84.0867
R1954 variable_delay_unit_8.forward.n2 variable_delay_unit_8.forward 19.8934
R1955 variable_delay_unit_8.forward variable_delay_unit_8.forward.n2 0.851271
R1956 variable_delay_unit_8.forward.n2 variable_delay_unit_8.forward.n1 0.465495
R1957 en_5.n0 en_5.t2 628.097
R1958 en_5.n1 en_5.t1 622.766
R1959 en_5.n2 en_5.t5 543.053
R1960 en_5.n0 en_5.t4 523.774
R1961 en_5.n4 en_5.t7 304.647
R1962 en_5.n4 en_5.t0 304.647
R1963 en_5.n2 en_5.t6 221.72
R1964 en_5 en_5.n2 220.304
R1965 en_5.n4 en_5.t3 202.44
R1966 en_5 en_5.n4 168.969
R1967 en_5 en_5.n1 166.147
R1968 en_5.n3 en_5 3.22371
R1969 en_5.n3 en_5 1.40175
R1970 en_5.n1 en_5.n0 1.09595
R1971 en_5 en_5.n3 0.443357
R1972 variable_delay_unit_2.in.n0 variable_delay_unit_2.in.t4 607.409
R1973 variable_delay_unit_2.in.n2 variable_delay_unit_2.in.t2 543.053
R1974 variable_delay_unit_2.in.n0 variable_delay_unit_2.in.t5 321.423
R1975 variable_delay_unit_2.in variable_delay_unit_2.in.n2 221.778
R1976 variable_delay_unit_2.in.n2 variable_delay_unit_2.in.t3 221.72
R1977 variable_delay_unit_2.in variable_delay_unit_2.in.n0 161.72
R1978 variable_delay_unit_2.in.n1 variable_delay_unit_2.in.t1 84.7227
R1979 variable_delay_unit_2.in.n1 variable_delay_unit_2.in.t0 84.0867
R1980 variable_delay_unit_2.in.n3 variable_delay_unit_2.in 20.0791
R1981 variable_delay_unit_2.in variable_delay_unit_2.in.n3 0.851271
R1982 variable_delay_unit_2.in.n3 variable_delay_unit_2.in.n1 0.465495
R1983 en_0.n2 en_0.t0 628.097
R1984 en_0.n3 en_0.t6 622.766
R1985 en_0.n0 en_0.t1 543.053
R1986 en_0.n2 en_0.t4 523.774
R1987 en_0.n1 en_0.t3 304.647
R1988 en_0.n1 en_0.t5 304.647
R1989 en_0.n0 en_0.t2 221.72
R1990 en_0.n5 en_0.n0 220.263
R1991 en_0.n1 en_0.t7 202.44
R1992 en_0 en_0.n1 168.969
R1993 en_0 en_0.n3 166.147
R1994 en_0 en_0.n4 3.17729
R1995 en_0.n4 en_0 1.40175
R1996 en_0.n3 en_0.n2 1.09595
R1997 en_0.n4 en_0 0.443357
R1998 en_0.n5 en_0 0.088
R1999 en_0 en_0.n5 0.063
R2000 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t6 628.097
R2001 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.t7 622.766
R2002 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t4 523.774
R2003 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t3 304.647
R2004 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t2 304.647
R2005 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t5 202.44
R2006 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n0 168.969
R2007 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n4 166.147
R2008 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t1 84.7557
R2009 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t0 84.1197
R2010 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R2011 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en 5.58443
R2012 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n2 4.59003
R2013 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.n3 1.09595
R2014 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t3 628.097
R2015 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.t5 622.766
R2016 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t7 523.774
R2017 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t6 304.647
R2018 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t2 304.647
R2019 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t4 202.44
R2020 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n0 168.969
R2021 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n4 166.147
R2022 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R2023 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R2024 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R2025 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en 5.58443
R2026 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n2 4.59003
R2027 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.n3 1.09595
R2028 en_4.n0 en_4.t2 628.097
R2029 en_4.n1 en_4.t0 622.766
R2030 en_4.n2 en_4.t5 543.053
R2031 en_4.n0 en_4.t4 523.774
R2032 en_4.n4 en_4.t3 304.647
R2033 en_4.n4 en_4.t7 304.647
R2034 en_4.n2 en_4.t6 221.72
R2035 en_4 en_4.n2 220.304
R2036 en_4.n4 en_4.t1 202.44
R2037 en_4 en_4.n4 168.969
R2038 en_4 en_4.n1 166.147
R2039 en_4.n3 en_4 3.22371
R2040 en_4.n3 en_4 1.40175
R2041 en_4.n1 en_4.n0 1.09595
R2042 en_4 en_4.n3 0.443357
R2043 variable_delay_unit_5.in.n0 variable_delay_unit_5.in.t4 607.409
R2044 variable_delay_unit_5.in.n2 variable_delay_unit_5.in.t2 543.053
R2045 variable_delay_unit_5.in.n0 variable_delay_unit_5.in.t5 321.423
R2046 variable_delay_unit_5.in variable_delay_unit_5.in.n2 221.778
R2047 variable_delay_unit_5.in.n2 variable_delay_unit_5.in.t3 221.72
R2048 variable_delay_unit_5.in variable_delay_unit_5.in.n0 161.72
R2049 variable_delay_unit_5.in.n1 variable_delay_unit_5.in.t1 84.7227
R2050 variable_delay_unit_5.in.n1 variable_delay_unit_5.in.t0 84.0867
R2051 variable_delay_unit_5.in.n3 variable_delay_unit_5.in 20.0791
R2052 variable_delay_unit_5.in variable_delay_unit_5.in.n3 0.851271
R2053 variable_delay_unit_5.in.n3 variable_delay_unit_5.in.n1 0.465495
R2054 variable_delay_unit_6.in.n0 variable_delay_unit_6.in.t4 607.409
R2055 variable_delay_unit_6.in.n2 variable_delay_unit_6.in.t2 543.053
R2056 variable_delay_unit_6.in.n0 variable_delay_unit_6.in.t5 321.423
R2057 variable_delay_unit_6.in variable_delay_unit_6.in.n2 221.778
R2058 variable_delay_unit_6.in.n2 variable_delay_unit_6.in.t3 221.72
R2059 variable_delay_unit_6.in variable_delay_unit_6.in.n0 161.72
R2060 variable_delay_unit_6.in.n1 variable_delay_unit_6.in.t1 84.7227
R2061 variable_delay_unit_6.in.n1 variable_delay_unit_6.in.t0 84.0867
R2062 variable_delay_unit_6.in.n3 variable_delay_unit_6.in 20.0791
R2063 variable_delay_unit_6.in variable_delay_unit_6.in.n3 0.851271
R2064 variable_delay_unit_6.in.n3 variable_delay_unit_6.in.n1 0.465495
R2065 en_3.n2 en_3.t0 628.097
R2066 en_3.n3 en_3.t7 622.766
R2067 en_3.n0 en_3.t3 543.053
R2068 en_3.n2 en_3.t2 523.774
R2069 en_3.n1 en_3.t5 304.647
R2070 en_3.n1 en_3.t6 304.647
R2071 en_3.n0 en_3.t4 221.72
R2072 en_3.n5 en_3.n0 220.263
R2073 en_3.n1 en_3.t1 202.44
R2074 en_3 en_3.n1 168.969
R2075 en_3 en_3.n3 166.147
R2076 en_3 en_3.n4 3.15229
R2077 en_3.n4 en_3 1.40175
R2078 en_3.n3 en_3.n2 1.09595
R2079 en_3.n4 en_3 0.443357
R2080 en_3.n5 en_3 0.113
R2081 en_3 en_3.n5 0.063
R2082 en_2.n2 en_2.t1 628.097
R2083 en_2.n3 en_2.t7 622.766
R2084 en_2.n0 en_2.t3 543.053
R2085 en_2.n2 en_2.t4 523.774
R2086 en_2.n1 en_2.t2 304.647
R2087 en_2.n1 en_2.t6 304.647
R2088 en_2.n0 en_2.t5 221.72
R2089 en_2.n5 en_2.n0 220.263
R2090 en_2.n1 en_2.t0 202.44
R2091 en_2 en_2.n1 168.969
R2092 en_2 en_2.n3 166.147
R2093 en_2 en_2.n4 3.09157
R2094 en_2.n4 en_2 1.40175
R2095 en_2.n3 en_2.n2 1.09595
R2096 en_2.n4 en_2 0.443357
R2097 en_2.n5 en_2 0.173714
R2098 en_2 en_2.n5 0.063
R2099 en_7.n0 en_7.t6 628.097
R2100 en_7.n1 en_7.t5 622.766
R2101 en_7.n2 en_7.t0 543.053
R2102 en_7.n0 en_7.t1 523.774
R2103 en_7.n4 en_7.t4 304.647
R2104 en_7.n4 en_7.t3 304.647
R2105 en_7.n2 en_7.t2 221.72
R2106 en_7 en_7.n2 220.304
R2107 en_7.n4 en_7.t7 202.44
R2108 en_7 en_7.n4 168.969
R2109 en_7 en_7.n1 166.147
R2110 en_7.n3 en_7 3.22371
R2111 en_7.n3 en_7 1.40175
R2112 en_7.n1 en_7.n0 1.09595
R2113 en_7 en_7.n3 0.443357
R2114 variable_delay_unit_7.tristate_inverter_1.en.n3 variable_delay_unit_7.tristate_inverter_1.en.t4 628.097
R2115 variable_delay_unit_7.tristate_inverter_1.en.n4 variable_delay_unit_7.tristate_inverter_1.en.t3 622.766
R2116 variable_delay_unit_7.tristate_inverter_1.en.n3 variable_delay_unit_7.tristate_inverter_1.en.t7 523.774
R2117 variable_delay_unit_7.tristate_inverter_1.en.n0 variable_delay_unit_7.tristate_inverter_1.en.t5 304.647
R2118 variable_delay_unit_7.tristate_inverter_1.en.n0 variable_delay_unit_7.tristate_inverter_1.en.t6 304.647
R2119 variable_delay_unit_7.tristate_inverter_1.en.n0 variable_delay_unit_7.tristate_inverter_1.en.t2 202.44
R2120 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_7.tristate_inverter_1.en.n0 168.969
R2121 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_7.tristate_inverter_1.en.n4 166.147
R2122 variable_delay_unit_7.tristate_inverter_1.en.n1 variable_delay_unit_7.tristate_inverter_1.en.t1 84.7557
R2123 variable_delay_unit_7.tristate_inverter_1.en.n1 variable_delay_unit_7.tristate_inverter_1.en.t0 84.1197
R2124 variable_delay_unit_7.tristate_inverter_1.en.n2 variable_delay_unit_7.tristate_inverter_1.en.n1 12.6535
R2125 variable_delay_unit_7.tristate_inverter_1.en.n2 variable_delay_unit_7.tristate_inverter_1.en 5.58443
R2126 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_7.tristate_inverter_1.en.n2 4.59003
R2127 variable_delay_unit_7.tristate_inverter_1.en.n4 variable_delay_unit_7.tristate_inverter_1.en.n3 1.09595
R2128 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t2 607.409
R2129 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t4 543.053
R2130 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t3 321.423
R2131 variable_delay_unit_1.in variable_delay_unit_1.in.n2 221.778
R2132 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t5 221.72
R2133 variable_delay_unit_1.in variable_delay_unit_1.in.n0 161.72
R2134 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t0 84.7227
R2135 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t1 84.0867
R2136 variable_delay_unit_1.in.n3 variable_delay_unit_1.in 20.0791
R2137 variable_delay_unit_1.in variable_delay_unit_1.in.n3 0.851271
R2138 variable_delay_unit_1.in.n3 variable_delay_unit_1.in.n1 0.465495
R2139 out.n0 out.t2 84.8477
R2140 out.n2 out.t0 84.8477
R2141 out.n0 out.t3 84.2063
R2142 out.n2 out.t1 84.1683
R2143 out out.n3 10.0241
R2144 out.n1 out 0.681535
R2145 out out.n0 0.287138
R2146 out.n3 out 0.0803611
R2147 out.n3 out.n2 0.0508472
R2148 out.n1 out 0.013431
R2149 out out.n1 0.0109167
R2150 variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_unit_4.tristate_inverter_1.en.t5 628.097
R2151 variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_unit_4.tristate_inverter_1.en.t7 622.766
R2152 variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_unit_4.tristate_inverter_1.en.t3 523.774
R2153 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t2 304.647
R2154 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t4 304.647
R2155 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t6 202.44
R2156 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n0 168.969
R2157 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n4 166.147
R2158 variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_unit_4.tristate_inverter_1.en.t1 84.7557
R2159 variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_unit_4.tristate_inverter_1.en.t0 84.1197
R2160 variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_unit_4.tristate_inverter_1.en.n1 12.6535
R2161 variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_unit_4.tristate_inverter_1.en 5.58443
R2162 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n2 4.59003
R2163 variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_unit_4.tristate_inverter_1.en.n3 1.09595
R2164 variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_unit_3.tristate_inverter_1.en.t5 628.097
R2165 variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_unit_3.tristate_inverter_1.en.t6 622.766
R2166 variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_unit_3.tristate_inverter_1.en.t3 523.774
R2167 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t7 304.647
R2168 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t2 304.647
R2169 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t4 202.44
R2170 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n0 168.969
R2171 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n4 166.147
R2172 variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_unit_3.tristate_inverter_1.en.t1 84.7557
R2173 variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_unit_3.tristate_inverter_1.en.t0 84.1197
R2174 variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_unit_3.tristate_inverter_1.en.n1 12.6535
R2175 variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_unit_3.tristate_inverter_1.en 5.58443
R2176 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n2 4.59003
R2177 variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_unit_3.tristate_inverter_1.en.n3 1.09595
R2178 variable_delay_unit_6.tristate_inverter_1.en.n3 variable_delay_unit_6.tristate_inverter_1.en.t5 628.097
R2179 variable_delay_unit_6.tristate_inverter_1.en.n4 variable_delay_unit_6.tristate_inverter_1.en.t7 622.766
R2180 variable_delay_unit_6.tristate_inverter_1.en.n3 variable_delay_unit_6.tristate_inverter_1.en.t3 523.774
R2181 variable_delay_unit_6.tristate_inverter_1.en.n0 variable_delay_unit_6.tristate_inverter_1.en.t4 304.647
R2182 variable_delay_unit_6.tristate_inverter_1.en.n0 variable_delay_unit_6.tristate_inverter_1.en.t6 304.647
R2183 variable_delay_unit_6.tristate_inverter_1.en.n0 variable_delay_unit_6.tristate_inverter_1.en.t2 202.44
R2184 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_6.tristate_inverter_1.en.n0 168.969
R2185 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_6.tristate_inverter_1.en.n4 166.147
R2186 variable_delay_unit_6.tristate_inverter_1.en.n1 variable_delay_unit_6.tristate_inverter_1.en.t1 84.7557
R2187 variable_delay_unit_6.tristate_inverter_1.en.n1 variable_delay_unit_6.tristate_inverter_1.en.t0 84.1197
R2188 variable_delay_unit_6.tristate_inverter_1.en.n2 variable_delay_unit_6.tristate_inverter_1.en.n1 12.6535
R2189 variable_delay_unit_6.tristate_inverter_1.en.n2 variable_delay_unit_6.tristate_inverter_1.en 5.58443
R2190 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_6.tristate_inverter_1.en.n2 4.59003
R2191 variable_delay_unit_6.tristate_inverter_1.en.n4 variable_delay_unit_6.tristate_inverter_1.en.n3 1.09595
R2192 variable_delay_unit_7.in.n0 variable_delay_unit_7.in.t2 607.409
R2193 variable_delay_unit_7.in.n2 variable_delay_unit_7.in.t3 543.053
R2194 variable_delay_unit_7.in.n0 variable_delay_unit_7.in.t4 321.423
R2195 variable_delay_unit_7.in variable_delay_unit_7.in.n2 221.778
R2196 variable_delay_unit_7.in.n2 variable_delay_unit_7.in.t5 221.72
R2197 variable_delay_unit_7.in variable_delay_unit_7.in.n0 161.72
R2198 variable_delay_unit_7.in.n1 variable_delay_unit_7.in.t1 84.7227
R2199 variable_delay_unit_7.in.n1 variable_delay_unit_7.in.t0 84.0867
R2200 variable_delay_unit_7.in.n3 variable_delay_unit_7.in 20.0791
R2201 variable_delay_unit_7.in variable_delay_unit_7.in.n3 0.851271
R2202 variable_delay_unit_7.in.n3 variable_delay_unit_7.in.n1 0.465495
R2203 in.n0 in.t0 543.053
R2204 in.n0 in.t1 221.72
R2205 in in.n0 221.565
R2206 variable_delay_unit_8.in.n0 variable_delay_unit_8.in.t3 607.409
R2207 variable_delay_unit_8.in.n2 variable_delay_unit_8.in.t2 543.053
R2208 variable_delay_unit_8.in.n0 variable_delay_unit_8.in.t5 321.423
R2209 variable_delay_unit_8.in variable_delay_unit_8.in.n2 221.778
R2210 variable_delay_unit_8.in.n2 variable_delay_unit_8.in.t4 221.72
R2211 variable_delay_unit_8.in variable_delay_unit_8.in.n0 161.72
R2212 variable_delay_unit_8.in.n1 variable_delay_unit_8.in.t1 84.7227
R2213 variable_delay_unit_8.in.n1 variable_delay_unit_8.in.t0 84.0867
R2214 variable_delay_unit_8.in.n3 variable_delay_unit_8.in 20.0791
R2215 variable_delay_unit_8.in variable_delay_unit_8.in.n3 0.851271
R2216 variable_delay_unit_8.in.n3 variable_delay_unit_8.in.n1 0.465495
C0 en_1 variable_delay_unit_2.tristate_inverter_1.en 1.5e-19
C1 variable_delay_unit_6.tristate_inverter_1.en a_19302_772# 0.11539f
C2 variable_delay_unit_2.in variable_delay_unit_1.in 0.087283f
C3 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.in 0.09141f
C4 a_5444_352# en_1 0.001909f
C5 a_2496_772# en_0 0.124274f
C6 variable_delay_unit_1.in in 0.08442f
C7 a_20184_772# variable_delay_unit_6.out 0.493816f
C8 VDD variable_delay_unit_4.in 2.12807f
C9 a_8392_352# en_2 0.001909f
C10 VDD a_20184_772# 1.6584f
C11 en_4 variable_delay_unit_3.out 2.67e-19
C12 a_23132_352# variable_delay_unit_8.out 0.070146f
C13 variable_delay_unit_8.out variable_delay_unit_8.tristate_inverter_1.en 0.12029f
C14 variable_delay_unit_5.out variable_delay_unit_4.tristate_inverter_1.en 0.085059f
C15 a_11340_772# a_11340_352# 0.011184f
C16 VDD variable_delay_unit_2.in 2.12807f
C17 a_14288_352# a_14288_772# 0.011184f
C18 a_10458_352# variable_delay_unit_4.in 0.054206f
C19 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_7.in 0.09141f
C20 VDD variable_delay_unit_1.tristate_inverter_1.en 2.77611f
C21 a_7510_352# variable_delay_unit_2.in 8.82e-20
C22 VDD in 0.238594f
C23 VDD variable_delay_unit_5.in 2.12807f
C24 variable_delay_unit_6.out a_20184_352# 0.172055f
C25 en_6 a_19302_772# 0.042718f
C26 VDD en_4 1.40792f
C27 VDD a_20184_352# 0.001468f
C28 en_1 a_4562_772# 0.042718f
C29 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.out 0.12029f
C30 variable_delay_unit_0.tristate_inverter_1.en a_2496_352# 0.15982f
C31 en_5 a_14288_352# 6.99e-20
C32 a_16354_352# en_5 0.15982f
C33 variable_delay_unit_6.in a_19302_772# 8.82e-20
C34 en_3 variable_delay_unit_3.out 0.224474f
C35 variable_delay_unit_0.tristate_inverter_1.en a_2496_772# 0.029284f
C36 variable_delay_unit_8.in variable_delay_unit_7.in 0.087283f
C37 a_23132_352# en_7 0.001909f
C38 variable_delay_unit_8.tristate_inverter_1.en a_25198_352# 2.39e-19
C39 variable_delay_unit_8.tristate_inverter_1.en en_7 1.5e-19
C40 a_17236_352# a_17236_772# 0.011184f
C41 a_16354_352# variable_delay_unit_5.tristate_inverter_1.en 2.39e-19
C42 a_23132_352# a_23132_772# 0.011184f
C43 a_13406_352# variable_delay_unit_4.out 0.222585f
C44 VDD en_3 1.40792f
C45 en_2 a_7510_772# 0.042718f
C46 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.in 0.09141f
C47 a_22250_772# en_7 0.042718f
C48 variable_delay_unit_8.forward a_26080_772# 0.016896f
C49 en_3 a_10458_352# 0.15982f
C50 a_5444_772# variable_delay_unit_2.out 0.071074f
C51 variable_delay_unit_3.out variable_delay_unit_4.out 0.071795f
C52 variable_delay_unit_3.in a_8392_772# 0.020173f
C53 variable_delay_unit_5.out variable_delay_unit_6.out 0.071795f
C54 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_8.forward 7.91e-21
C55 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C56 VDD variable_delay_unit_5.out 1.34424f
C57 variable_delay_unit_3.in variable_delay_unit_2.out 0.235667f
C58 a_16354_352# a_16354_772# 0.004142f
C59 a_16354_352# variable_delay_unit_6.in 0.054206f
C60 variable_delay_unit_3.in a_10458_772# 8.82e-20
C61 variable_delay_unit_6.out variable_delay_unit_7.out 0.071795f
C62 en_1 variable_delay_unit_2.out 0.043504f
C63 VDD variable_delay_unit_7.out 1.3445f
C64 VDD variable_delay_unit_4.out 1.34424f
C65 out a_2496_352# 0.172055f
C66 variable_delay_unit_4.in variable_delay_unit_5.in 0.087283f
C67 a_20184_772# a_20184_352# 0.011184f
C68 en_4 variable_delay_unit_4.in 0.506369f
C69 a_8392_772# variable_delay_unit_2.tristate_inverter_1.en 0.029284f
C70 a_22250_352# VDD 6.98e-19
C71 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.out 0.12029f
C72 a_2496_772# out 0.493816f
C73 variable_delay_unit_8.forward variable_delay_unit_8.in 0.087283f
C74 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_2.in 0.814958f
C75 variable_delay_unit_1.out en_2 2.67e-19
C76 variable_delay_unit_8.out a_26080_352# 0.172055f
C77 a_5444_352# variable_delay_unit_2.out 0.070146f
C78 en_5 a_17236_352# 0.001909f
C79 en_4 variable_delay_unit_5.in 0.574722f
C80 en_2 variable_delay_unit_3.out 0.043504f
C81 en_1 en_0 0.010459f
C82 a_14288_772# variable_delay_unit_4.tristate_inverter_1.en 0.029284f
C83 variable_delay_unit_8.tristate_inverter_1.en a_26080_772# 0.029284f
C84 variable_delay_unit_5.tristate_inverter_1.en a_17236_352# 0.15982f
C85 en_3 variable_delay_unit_4.in 0.574722f
C86 a_11340_352# variable_delay_unit_3.in 7.65e-21
C87 a_23132_352# variable_delay_unit_7.tristate_inverter_1.en 0.15982f
C88 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_8.tristate_inverter_1.en 0.002365f
C89 en_5 variable_delay_unit_4.tristate_inverter_1.en 9.38e-20
C90 variable_delay_unit_8.out a_25198_772# 0.505512f
C91 VDD en_2 1.40792f
C92 a_17236_772# variable_delay_unit_6.out 0.071074f
C93 a_7510_352# en_2 0.15982f
C94 VDD a_17236_772# 1.6584f
C95 variable_delay_unit_7.in a_19302_772# 0.088132f
C96 en_3 variable_delay_unit_5.in 3.37e-20
C97 en_6 a_17236_352# 6.99e-20
C98 variable_delay_unit_1.out a_2496_352# 0.070146f
C99 en_4 en_3 0.010459f
C100 variable_delay_unit_7.tristate_inverter_1.en a_22250_772# 0.11539f
C101 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en 0.002365f
C102 a_2496_772# variable_delay_unit_1.out 0.071074f
C103 variable_delay_unit_0.tristate_inverter_1.en en_1 9.38e-20
C104 variable_delay_unit_8.in variable_delay_unit_8.tristate_inverter_1.en 0.09141f
C105 a_20184_772# variable_delay_unit_7.out 0.071074f
C106 a_11340_772# variable_delay_unit_3.out 0.493816f
C107 VDD variable_delay_unit_8.out 1.5668f
C108 variable_delay_unit_4.in variable_delay_unit_4.out 0.499092f
C109 a_2496_772# variable_delay_unit_1.in 0.020173f
C110 variable_delay_unit_5.out variable_delay_unit_5.in 0.499092f
C111 en_0 a_1614_352# 0.15982f
C112 en_4 variable_delay_unit_5.out 0.043504f
C113 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_2.out 0.002141f
C114 variable_delay_unit_8.in a_22250_772# 0.088132f
C115 a_25198_352# a_25198_772# 0.004142f
C116 VDD a_2496_352# 0.001468f
C117 variable_delay_unit_3.tristate_inverter_1.en a_10458_772# 0.11539f
C118 a_20184_352# variable_delay_unit_7.out 0.070146f
C119 a_11340_772# VDD 1.6584f
C120 variable_delay_unit_5.in variable_delay_unit_4.out 0.235667f
C121 en_4 variable_delay_unit_4.out 0.224474f
C122 VDD a_2496_772# 1.6584f
C123 a_8392_352# variable_delay_unit_2.tristate_inverter_1.en 0.15982f
C124 variable_delay_unit_6.in variable_delay_unit_4.tristate_inverter_1.en 7.91e-21
C125 VDD a_14288_772# 1.6584f
C126 a_8392_772# variable_delay_unit_2.out 0.493816f
C127 variable_delay_unit_6.out en_7 2.67e-19
C128 VDD a_25198_352# 0.160518f
C129 VDD en_7 1.41838f
C130 en_5 variable_delay_unit_6.out 0.043504f
C131 a_23132_352# variable_delay_unit_7.in 7.65e-21
C132 VDD en_5 1.40792f
C133 variable_delay_unit_0.tristate_inverter_1.en a_1614_352# 2.39e-19
C134 VDD a_23132_772# 1.65847f
C135 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_6.out 0.12029f
C136 VDD variable_delay_unit_6.tristate_inverter_1.en 2.77611f
C137 variable_delay_unit_4.in en_2 3.37e-20
C138 a_7510_772# variable_delay_unit_3.in 0.088132f
C139 en_3 variable_delay_unit_4.out 0.043504f
C140 variable_delay_unit_7.in a_22250_772# 8.82e-20
C141 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_6.out 0.085059f
C142 VDD variable_delay_unit_5.tristate_inverter_1.en 2.77611f
C143 en_1 out 2.67e-19
C144 a_26080_352# a_26080_772# 0.011184f
C145 variable_delay_unit_2.in en_2 0.506369f
C146 variable_delay_unit_1.tristate_inverter_1.en en_2 9.38e-20
C147 en_1 a_4562_352# 0.15982f
C148 variable_delay_unit_3.tristate_inverter_1.en a_11340_352# 0.15982f
C149 a_17236_772# variable_delay_unit_5.in 7.65e-21
C150 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en 0.11539f
C151 en_6 variable_delay_unit_6.out 0.224474f
C152 VDD en_6 1.40792f
C153 variable_delay_unit_5.out variable_delay_unit_4.out 0.071795f
C154 variable_delay_unit_6.tristate_inverter_1.en a_19302_352# 2.39e-19
C155 variable_delay_unit_6.in variable_delay_unit_6.out 0.499092f
C156 a_11340_772# variable_delay_unit_4.in 0.020173f
C157 VDD a_16354_772# 1.6584f
C158 VDD variable_delay_unit_6.in 2.12807f
C159 a_22250_352# variable_delay_unit_7.out 0.222585f
C160 variable_delay_unit_8.in a_26080_352# 7.65e-21
C161 en_3 en_2 0.010459f
C162 a_1614_772# a_1614_352# 0.004142f
C163 variable_delay_unit_1.out a_5444_772# 0.493816f
C164 variable_delay_unit_8.forward variable_delay_unit_8.tristate_inverter_1.en 0.794183f
C165 a_14288_772# variable_delay_unit_4.in 7.65e-21
C166 in a_2496_352# 7.65e-21
C167 a_4562_352# a_4562_772# 0.004142f
C168 out a_1614_352# 0.222585f
C169 en_6 a_19302_352# 0.15982f
C170 a_11340_772# en_4 6.99e-20
C171 variable_delay_unit_1.in a_5444_772# 7.65e-21
C172 a_2496_772# in 7.65e-21
C173 en_1 variable_delay_unit_1.out 0.224474f
C174 a_20184_772# en_7 6.99e-20
C175 VDD a_26080_772# 1.78268f
C176 a_8392_352# a_8392_772# 0.011184f
C177 a_14288_772# variable_delay_unit_5.in 0.020173f
C178 variable_delay_unit_3.out variable_delay_unit_3.in 0.499092f
C179 en_4 a_14288_772# 0.124274f
C180 a_8392_352# variable_delay_unit_2.out 0.172055f
C181 a_20184_772# variable_delay_unit_6.tristate_inverter_1.en 0.029284f
C182 en_1 variable_delay_unit_1.in 0.506369f
C183 variable_delay_unit_8.in a_25198_772# 8.82e-20
C184 variable_delay_unit_6.in a_19302_352# 8.82e-20
C185 variable_delay_unit_1.out variable_delay_unit_2.tristate_inverter_1.en 0.002141f
C186 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_6.out 0.002141f
C187 a_17236_772# variable_delay_unit_5.out 0.493816f
C188 VDD variable_delay_unit_7.tristate_inverter_1.en 2.7762f
C189 VDD a_5444_772# 1.6584f
C190 en_5 variable_delay_unit_5.in 0.506369f
C191 a_20184_352# en_7 6.99e-20
C192 en_4 en_5 0.010459f
C193 a_5444_352# variable_delay_unit_1.out 0.172055f
C194 VDD variable_delay_unit_3.in 2.12807f
C195 variable_delay_unit_0.tristate_inverter_1.en en_0 1.09349f
C196 a_7510_352# variable_delay_unit_3.in 0.054206f
C197 variable_delay_unit_3.out variable_delay_unit_2.tristate_inverter_1.en 0.085059f
C198 variable_delay_unit_6.tristate_inverter_1.en a_20184_352# 0.15982f
C199 a_11340_772# en_3 0.124274f
C200 VDD en_1 1.40792f
C201 a_5444_352# variable_delay_unit_1.in 7.65e-21
C202 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.in 0.09141f
C203 a_10458_352# variable_delay_unit_3.in 8.82e-20
C204 en_4 variable_delay_unit_5.tristate_inverter_1.en 1.5e-19
C205 VDD variable_delay_unit_8.in 2.63444f
C206 a_20184_772# en_6 0.124274f
C207 VDD variable_delay_unit_2.tristate_inverter_1.en 2.77611f
C208 variable_delay_unit_1.out a_4562_772# 0.505512f
C209 variable_delay_unit_8.out variable_delay_unit_7.out 0.071795f
C210 a_7510_352# variable_delay_unit_2.tristate_inverter_1.en 2.39e-19
C211 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en 0.002365f
C212 VDD a_5444_352# 0.001468f
C213 a_20184_772# variable_delay_unit_6.in 7.65e-21
C214 variable_delay_unit_1.in a_4562_772# 8.82e-20
C215 en_6 a_20184_352# 0.001909f
C216 a_7510_772# variable_delay_unit_2.out 0.505512f
C217 variable_delay_unit_1.in a_1614_352# 0.054206f
C218 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en 0.11539f
C219 variable_delay_unit_5.out a_14288_772# 0.071074f
C220 a_11340_772# variable_delay_unit_4.out 0.071074f
C221 a_16354_772# variable_delay_unit_5.in 8.82e-20
C222 variable_delay_unit_6.in variable_delay_unit_5.in 0.087283f
C223 variable_delay_unit_6.in a_20184_352# 7.65e-21
C224 en_4 variable_delay_unit_6.in 3.37e-20
C225 VDD a_4562_772# 1.6584f
C226 a_14288_772# variable_delay_unit_4.out 0.493816f
C227 en_5 variable_delay_unit_5.out 0.224474f
C228 a_1614_772# en_0 0.042718f
C229 VDD a_1614_352# 6.98e-19
C230 variable_delay_unit_7.in variable_delay_unit_6.out 0.235667f
C231 en_7 variable_delay_unit_7.out 0.224474f
C232 VDD variable_delay_unit_7.in 2.12807f
C233 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_5.out 0.002141f
C234 en_0 out 0.218964f
C235 en_5 variable_delay_unit_4.out 2.67e-19
C236 variable_delay_unit_7.out a_23132_772# 0.493816f
C237 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_7.out 0.085059f
C238 a_13406_352# a_13406_772# 0.004142f
C239 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.out 0.12029f
C240 a_22250_352# en_7 0.15982f
C241 variable_delay_unit_4.in variable_delay_unit_3.in 0.087283f
C242 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.out 0.12029f
C243 variable_delay_unit_2.in a_5444_772# 0.020173f
C244 variable_delay_unit_1.tristate_inverter_1.en a_5444_772# 0.029284f
C245 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_4.out 0.002141f
C246 variable_delay_unit_1.out variable_delay_unit_2.out 0.071795f
C247 variable_delay_unit_2.in variable_delay_unit_3.in 0.087283f
C248 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_3.in 7.91e-21
C249 en_6 variable_delay_unit_5.out 2.67e-19
C250 a_14288_352# variable_delay_unit_4.tristate_inverter_1.en 0.15982f
C251 en_1 variable_delay_unit_2.in 0.574722f
C252 VDD variable_delay_unit_3.tristate_inverter_1.en 2.77611f
C253 variable_delay_unit_0.tristate_inverter_1.en a_1614_772# 0.11539f
C254 variable_delay_unit_7.in a_19302_352# 0.054206f
C255 variable_delay_unit_8.forward a_25198_772# 0.088132f
C256 en_1 variable_delay_unit_1.tristate_inverter_1.en 1.09349f
C257 variable_delay_unit_3.out a_8392_772# 0.071074f
C258 variable_delay_unit_4.in variable_delay_unit_2.tristate_inverter_1.en 7.91e-21
C259 variable_delay_unit_3.out variable_delay_unit_2.out 0.071795f
C260 en_6 variable_delay_unit_7.out 0.043504f
C261 variable_delay_unit_3.out a_10458_772# 0.505512f
C262 variable_delay_unit_0.tristate_inverter_1.en out 0.12022f
C263 variable_delay_unit_3.tristate_inverter_1.en a_10458_352# 2.39e-19
C264 variable_delay_unit_5.out a_16354_772# 0.505512f
C265 variable_delay_unit_2.in variable_delay_unit_2.tristate_inverter_1.en 0.09141f
C266 variable_delay_unit_6.in variable_delay_unit_5.out 0.235667f
C267 VDD a_13406_772# 1.6584f
C268 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C269 VDD a_8392_772# 1.6584f
C270 variable_delay_unit_6.out a_19302_772# 0.505512f
C271 VDD a_19302_772# 1.6584f
C272 en_5 a_17236_772# 0.124274f
C273 VDD variable_delay_unit_2.out 1.34424f
C274 a_5444_352# variable_delay_unit_1.tristate_inverter_1.en 0.15982f
C275 a_7510_352# variable_delay_unit_2.out 0.222585f
C276 variable_delay_unit_1.out en_0 0.043504f
C277 VDD a_10458_772# 1.6584f
C278 VDD variable_delay_unit_8.forward 2.28561f
C279 variable_delay_unit_8.tristate_inverter_1.en a_26080_352# 0.15982f
C280 en_3 variable_delay_unit_3.in 0.506369f
C281 variable_delay_unit_1.in en_0 0.574722f
C282 variable_delay_unit_5.tristate_inverter_1.en a_17236_772# 0.029284f
C283 a_10458_352# a_10458_772# 0.004142f
C284 a_2496_772# a_2496_352# 0.011184f
C285 variable_delay_unit_8.out a_25198_352# 0.222585f
C286 a_20184_772# variable_delay_unit_7.in 0.020173f
C287 variable_delay_unit_8.out en_7 0.043504f
C288 variable_delay_unit_2.in a_4562_772# 0.088132f
C289 variable_delay_unit_1.tristate_inverter_1.en a_4562_772# 0.11539f
C290 variable_delay_unit_8.out a_23132_772# 0.071074f
C291 en_3 variable_delay_unit_2.tristate_inverter_1.en 9.38e-20
C292 in a_1614_352# 8.82e-20
C293 a_19302_772# a_19302_352# 0.004142f
C294 VDD en_0 1.41013f
C295 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_7.out 0.12029f
C296 variable_delay_unit_8.tristate_inverter_1.en a_25198_772# 0.11539f
C297 en_6 a_17236_772# 6.99e-20
C298 a_11340_352# variable_delay_unit_3.out 0.172055f
C299 a_1614_772# out 0.505512f
C300 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.out 0.085059f
C301 VDD a_14288_352# 0.001468f
C302 VDD a_16354_352# 6.98e-19
C303 a_22250_352# variable_delay_unit_7.tristate_inverter_1.en 2.39e-19
C304 en_5 a_14288_772# 6.99e-20
C305 variable_delay_unit_6.in a_17236_772# 0.020173f
C306 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.in 0.814958f
C307 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.in 0.814958f
C308 VDD a_11340_352# 0.001468f
C309 variable_delay_unit_8.in variable_delay_unit_7.out 0.235667f
C310 a_23132_352# VDD 0.001538f
C311 VDD variable_delay_unit_8.tristate_inverter_1.en 3.86957f
C312 a_13406_772# variable_delay_unit_4.in 8.82e-20
C313 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_5.in 7.91e-21
C314 en_7 a_23132_772# 0.124274f
C315 variable_delay_unit_6.tristate_inverter_1.en en_7 9.38e-20
C316 a_8392_352# variable_delay_unit_3.out 0.070146f
C317 en_4 variable_delay_unit_3.tristate_inverter_1.en 9.38e-20
C318 a_22250_352# variable_delay_unit_8.in 0.054206f
C319 VDD variable_delay_unit_0.tristate_inverter_1.en 2.77513f
C320 en_5 variable_delay_unit_6.tristate_inverter_1.en 1.5e-19
C321 VDD a_22250_772# 1.6584f
C322 variable_delay_unit_4.in a_10458_772# 0.088132f
C323 en_5 variable_delay_unit_5.tristate_inverter_1.en 1.09349f
C324 a_13406_772# variable_delay_unit_5.in 0.088132f
C325 variable_delay_unit_2.in a_8392_772# 7.65e-21
C326 en_2 a_5444_772# 6.99e-20
C327 en_4 a_13406_772# 0.042718f
C328 variable_delay_unit_2.in variable_delay_unit_2.out 0.499092f
C329 VDD a_8392_352# 0.001468f
C330 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_2.out 0.085059f
C331 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en 0.002365f
C332 en_2 variable_delay_unit_3.in 0.574722f
C333 en_6 en_7 0.010459f
C334 variable_delay_unit_8.out a_26080_772# 0.493816f
C335 en_1 en_2 0.010459f
C336 en_5 en_6 0.010459f
C337 variable_delay_unit_3.tristate_inverter_1.en en_3 1.09349f
C338 variable_delay_unit_7.in variable_delay_unit_7.out 0.499092f
C339 variable_delay_unit_1.out out 0.071795f
C340 variable_delay_unit_1.in a_1614_772# 0.088132f
C341 en_6 variable_delay_unit_6.tristate_inverter_1.en 1.09349f
C342 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_8.out 0.085059f
C343 variable_delay_unit_1.out a_4562_352# 0.222585f
C344 en_2 variable_delay_unit_2.tristate_inverter_1.en 1.09349f
C345 a_13406_352# variable_delay_unit_4.tristate_inverter_1.en 2.39e-19
C346 en_5 a_16354_772# 0.042718f
C347 a_22250_352# variable_delay_unit_7.in 8.82e-20
C348 en_5 variable_delay_unit_6.in 0.574722f
C349 variable_delay_unit_1.in out 0.235655f
C350 en_6 variable_delay_unit_5.tristate_inverter_1.en 9.38e-20
C351 variable_delay_unit_2.in en_0 3.37e-20
C352 a_14288_352# variable_delay_unit_4.in 7.65e-21
C353 a_5444_352# en_2 6.99e-20
C354 en_3 a_8392_772# 6.99e-20
C355 variable_delay_unit_1.in a_4562_352# 8.82e-20
C356 variable_delay_unit_1.tristate_inverter_1.en en_0 1.5e-19
C357 en_0 in 0.259572f
C358 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_6.in 0.09141f
C359 a_17236_352# variable_delay_unit_6.out 0.070146f
C360 VDD a_17236_352# 0.001468f
C361 en_3 variable_delay_unit_2.out 2.67e-19
C362 VDD a_1614_772# 1.6584f
C363 en_3 a_10458_772# 0.042718f
C364 variable_delay_unit_5.tristate_inverter_1.en a_16354_772# 0.11539f
C365 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_6.in 0.814958f
C366 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_3.out 0.002141f
C367 VDD out 1.15938f
C368 a_11340_772# variable_delay_unit_3.in 7.65e-21
C369 variable_delay_unit_8.in variable_delay_unit_8.out 0.499092f
C370 a_16354_352# variable_delay_unit_5.in 8.82e-20
C371 VDD a_7510_772# 1.6584f
C372 en_1 a_2496_352# 6.99e-20
C373 en_4 a_14288_352# 0.001909f
C374 a_7510_352# a_7510_772# 0.004142f
C375 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.out 0.085059f
C376 VDD a_4562_352# 6.98e-19
C377 en_4 a_11340_352# 6.99e-20
C378 en_1 a_2496_772# 6.99e-20
C379 variable_delay_unit_7.tristate_inverter_1.en en_7 1.09349f
C380 VDD variable_delay_unit_4.tristate_inverter_1.en 2.77611f
C381 en_6 variable_delay_unit_6.in 0.506369f
C382 a_13406_772# variable_delay_unit_4.out 0.505512f
C383 variable_delay_unit_7.tristate_inverter_1.en a_23132_772# 0.029284f
C384 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_2.in 7.91e-21
C385 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_7.tristate_inverter_1.en 0.002365f
C386 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en 0.002365f
C387 variable_delay_unit_0.tristate_inverter_1.en in 0.091118f
C388 VDD a_26080_352# 0.003377f
C389 variable_delay_unit_6.in a_16354_772# 0.088132f
C390 variable_delay_unit_1.in variable_delay_unit_1.out 0.499092f
C391 variable_delay_unit_8.in a_25198_352# 8.82e-20
C392 a_8392_352# variable_delay_unit_2.in 7.65e-21
C393 variable_delay_unit_8.in en_7 0.574722f
C394 a_11340_352# en_3 0.001909f
C395 VDD a_13406_352# 6.98e-19
C396 variable_delay_unit_8.in a_23132_772# 0.020173f
C397 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_8.in 7.91e-21
C398 variable_delay_unit_3.tristate_inverter_1.en en_2 1.5e-19
C399 en_6 variable_delay_unit_7.tristate_inverter_1.en 1.5e-19
C400 VDD variable_delay_unit_1.out 1.34424f
C401 VDD a_25198_772# 1.70112f
C402 a_14288_352# variable_delay_unit_5.out 0.070146f
C403 a_16354_352# variable_delay_unit_5.out 0.222585f
C404 VDD variable_delay_unit_1.in 2.12798f
C405 VDD variable_delay_unit_3.out 1.34424f
C406 en_2 a_8392_772# 0.124274f
C407 en_2 variable_delay_unit_2.out 0.224474f
C408 a_14288_352# variable_delay_unit_4.out 0.172055f
C409 en_3 a_8392_352# 6.99e-20
C410 en_6 variable_delay_unit_8.in 3.37e-20
C411 a_10458_352# variable_delay_unit_3.out 0.222585f
C412 a_1614_772# in 8.82e-20
C413 a_17236_352# variable_delay_unit_5.in 7.65e-21
C414 a_11340_352# variable_delay_unit_4.out 0.070146f
C415 VDD variable_delay_unit_6.out 1.34424f
C416 variable_delay_unit_7.in en_7 0.506369f
C417 en_5 variable_delay_unit_7.in 3.37e-20
C418 a_23132_352# variable_delay_unit_7.out 0.172055f
C419 variable_delay_unit_8.tristate_inverter_1.en variable_delay_unit_7.out 0.002141f
C420 a_7510_352# VDD 6.98e-19
C421 variable_delay_unit_1.tristate_inverter_1.en out 0.002141f
C422 variable_delay_unit_2.in a_7510_772# 8.82e-20
C423 in out 0.487038f
C424 variable_delay_unit_7.in a_23132_772# 7.65e-21
C425 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.in 0.09141f
C426 variable_delay_unit_2.in a_4562_352# 0.054206f
C427 variable_delay_unit_6.tristate_inverter_1.en variable_delay_unit_7.in 0.814958f
C428 variable_delay_unit_1.tristate_inverter_1.en a_4562_352# 2.39e-19
C429 a_11340_772# variable_delay_unit_3.tristate_inverter_1.en 0.029284f
C430 VDD a_10458_352# 6.98e-19
C431 a_22250_772# variable_delay_unit_7.out 0.505512f
C432 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_7.in 7.91e-21
C433 variable_delay_unit_8.forward variable_delay_unit_8.out 0.234428f
C434 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_5.in 0.814958f
C435 en_4 variable_delay_unit_4.tristate_inverter_1.en 1.09349f
C436 a_22250_352# a_22250_772# 0.004142f
C437 variable_delay_unit_8.in a_26080_772# 7.65e-21
C438 variable_delay_unit_6.out a_19302_352# 0.222585f
C439 VDD a_19302_352# 6.98e-19
C440 en_1 a_5444_772# 0.124274f
C441 a_13406_352# variable_delay_unit_4.in 8.82e-20
C442 en_6 variable_delay_unit_7.in 0.574722f
C443 en_1 variable_delay_unit_3.in 3.37e-20
C444 variable_delay_unit_7.tristate_inverter_1.en variable_delay_unit_8.in 0.814958f
C445 variable_delay_unit_6.in variable_delay_unit_7.in 0.087283f
C446 a_13406_352# variable_delay_unit_5.in 0.054206f
C447 variable_delay_unit_3.in variable_delay_unit_2.tristate_inverter_1.en 0.814958f
C448 en_4 a_13406_352# 0.15982f
C449 a_17236_352# variable_delay_unit_5.out 0.172055f
C450 a_5444_352# a_5444_772# 0.011184f
C451 variable_delay_unit_2.in variable_delay_unit_1.out 0.235667f
C452 en_3 variable_delay_unit_4.tristate_inverter_1.en 1.5e-19
C453 variable_delay_unit_4.in variable_delay_unit_3.out 0.235667f
C454 variable_delay_unit_8.forward a_25198_352# 0.054206f
C455 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.out 0.12029f
C456 variable_delay_unit_8.forward en_7 3.37e-20
C457 en_0 a_2496_352# 0.001909f
C458 en_7 VSS 2.08969f
C459 en_6 VSS 2.08969f
C460 en_5 VSS 2.08969f
C461 en_4 VSS 2.08969f
C462 en_3 VSS 2.08969f
C463 en_2 VSS 2.08969f
C464 en_1 VSS 2.08969f
C465 out VSS 1.89289f
C466 in VSS 1.0591f
C467 en_0 VSS 2.22578f
C468 VDD VSS 77.568855f
C469 a_26080_352# VSS 0.783967f
C470 a_25198_352# VSS 0.71648f
C471 a_23132_352# VSS 0.717347f
C472 a_22250_352# VSS 0.71648f
C473 a_26080_772# VSS 0.114203f
C474 a_25198_772# VSS 0.037888f
C475 variable_delay_unit_8.forward VSS 2.632682f
C476 variable_delay_unit_8.tristate_inverter_1.en VSS 2.962211f
C477 a_20184_352# VSS 0.717347f
C478 a_19302_352# VSS 0.71648f
C479 a_23132_772# VSS 0.043128f
C480 variable_delay_unit_8.out VSS 2.29731f
C481 a_22250_772# VSS 0.037888f
C482 variable_delay_unit_8.in VSS 3.857309f
C483 variable_delay_unit_7.tristate_inverter_1.en VSS 2.51692f
C484 a_17236_352# VSS 0.717347f
C485 a_16354_352# VSS 0.71648f
C486 a_20184_772# VSS 0.043128f
C487 variable_delay_unit_7.out VSS 2.21957f
C488 a_19302_772# VSS 0.037888f
C489 variable_delay_unit_7.in VSS 3.60152f
C490 variable_delay_unit_6.tristate_inverter_1.en VSS 2.51692f
C491 a_14288_352# VSS 0.717347f
C492 a_13406_352# VSS 0.71648f
C493 a_17236_772# VSS 0.043128f
C494 variable_delay_unit_6.out VSS 2.21957f
C495 a_16354_772# VSS 0.037888f
C496 variable_delay_unit_6.in VSS 3.60152f
C497 variable_delay_unit_5.tristate_inverter_1.en VSS 2.51692f
C498 a_11340_352# VSS 0.717347f
C499 a_10458_352# VSS 0.71648f
C500 a_14288_772# VSS 0.043128f
C501 variable_delay_unit_5.out VSS 2.21957f
C502 a_13406_772# VSS 0.037888f
C503 variable_delay_unit_5.in VSS 3.60152f
C504 variable_delay_unit_4.tristate_inverter_1.en VSS 2.51692f
C505 a_8392_352# VSS 0.717347f
C506 a_7510_352# VSS 0.71648f
C507 a_11340_772# VSS 0.043128f
C508 variable_delay_unit_4.out VSS 2.21957f
C509 a_10458_772# VSS 0.037888f
C510 variable_delay_unit_4.in VSS 3.60152f
C511 variable_delay_unit_3.tristate_inverter_1.en VSS 2.51692f
C512 a_5444_352# VSS 0.717347f
C513 a_4562_352# VSS 0.71648f
C514 a_8392_772# VSS 0.043128f
C515 variable_delay_unit_3.out VSS 2.21957f
C516 a_7510_772# VSS 0.037888f
C517 variable_delay_unit_3.in VSS 3.60152f
C518 variable_delay_unit_2.tristate_inverter_1.en VSS 2.51692f
C519 a_2496_352# VSS 0.717347f
C520 a_1614_352# VSS 0.71648f
C521 a_5444_772# VSS 0.043128f
C522 variable_delay_unit_2.out VSS 2.21957f
C523 a_4562_772# VSS 0.037888f
C524 variable_delay_unit_2.in VSS 3.60152f
C525 variable_delay_unit_1.tristate_inverter_1.en VSS 2.51692f
C526 a_2496_772# VSS 0.043128f
C527 variable_delay_unit_1.out VSS 2.21957f
C528 a_1614_772# VSS 0.037888f
C529 variable_delay_unit_1.in VSS 3.60479f
C530 variable_delay_unit_0.tristate_inverter_1.en VSS 2.52279f
C531 variable_delay_unit_8.in.t3 VSS 0.055694f
C532 variable_delay_unit_8.in.t5 VSS 0.021119f
C533 variable_delay_unit_8.in.n0 VSS 0.058574f
C534 variable_delay_unit_8.in.t0 VSS 0.041029f
C535 variable_delay_unit_8.in.t1 VSS 0.130438f
C536 variable_delay_unit_8.in.n1 VSS 0.316137f
C537 variable_delay_unit_8.in.t2 VSS 0.053167f
C538 variable_delay_unit_8.in.t4 VSS 0.017162f
C539 variable_delay_unit_8.in.n2 VSS 0.055911f
C540 variable_delay_unit_8.in.n3 VSS 0.520657f
C541 variable_delay_unit_7.in.t2 VSS 0.044984f
C542 variable_delay_unit_7.in.t4 VSS 0.017058f
C543 variable_delay_unit_7.in.n0 VSS 0.04731f
C544 variable_delay_unit_7.in.t0 VSS 0.033139f
C545 variable_delay_unit_7.in.t1 VSS 0.105354f
C546 variable_delay_unit_7.in.n1 VSS 0.255341f
C547 variable_delay_unit_7.in.t3 VSS 0.042943f
C548 variable_delay_unit_7.in.t5 VSS 0.013862f
C549 variable_delay_unit_7.in.n2 VSS 0.045159f
C550 variable_delay_unit_7.in.n3 VSS 0.420531f
C551 variable_delay_unit_6.tristate_inverter_1.en.t2 VSS 0.019446f
C552 variable_delay_unit_6.tristate_inverter_1.en.t6 VSS 0.025128f
C553 variable_delay_unit_6.tristate_inverter_1.en.t4 VSS 0.025128f
C554 variable_delay_unit_6.tristate_inverter_1.en.n0 VSS 0.074066f
C555 variable_delay_unit_6.tristate_inverter_1.en.t1 VSS 0.154367f
C556 variable_delay_unit_6.tristate_inverter_1.en.t0 VSS 0.048564f
C557 variable_delay_unit_6.tristate_inverter_1.en.n1 VSS 0.616703f
C558 variable_delay_unit_6.tristate_inverter_1.en.n2 VSS 0.678061f
C559 variable_delay_unit_6.tristate_inverter_1.en.t7 VSS 0.066961f
C560 variable_delay_unit_6.tristate_inverter_1.en.t3 VSS 0.062029f
C561 variable_delay_unit_6.tristate_inverter_1.en.t5 VSS 0.067187f
C562 variable_delay_unit_6.tristate_inverter_1.en.n3 VSS 0.065756f
C563 variable_delay_unit_6.tristate_inverter_1.en.n4 VSS 0.045654f
C564 variable_delay_unit_3.tristate_inverter_1.en.t4 VSS 0.019446f
C565 variable_delay_unit_3.tristate_inverter_1.en.t2 VSS 0.025128f
C566 variable_delay_unit_3.tristate_inverter_1.en.t7 VSS 0.025128f
C567 variable_delay_unit_3.tristate_inverter_1.en.n0 VSS 0.074066f
C568 variable_delay_unit_3.tristate_inverter_1.en.t1 VSS 0.154367f
C569 variable_delay_unit_3.tristate_inverter_1.en.t0 VSS 0.048564f
C570 variable_delay_unit_3.tristate_inverter_1.en.n1 VSS 0.616703f
C571 variable_delay_unit_3.tristate_inverter_1.en.n2 VSS 0.678061f
C572 variable_delay_unit_3.tristate_inverter_1.en.t6 VSS 0.066961f
C573 variable_delay_unit_3.tristate_inverter_1.en.t3 VSS 0.062029f
C574 variable_delay_unit_3.tristate_inverter_1.en.t5 VSS 0.067187f
C575 variable_delay_unit_3.tristate_inverter_1.en.n3 VSS 0.065756f
C576 variable_delay_unit_3.tristate_inverter_1.en.n4 VSS 0.045654f
C577 variable_delay_unit_4.tristate_inverter_1.en.t6 VSS 0.019446f
C578 variable_delay_unit_4.tristate_inverter_1.en.t4 VSS 0.025128f
C579 variable_delay_unit_4.tristate_inverter_1.en.t2 VSS 0.025128f
C580 variable_delay_unit_4.tristate_inverter_1.en.n0 VSS 0.074066f
C581 variable_delay_unit_4.tristate_inverter_1.en.t1 VSS 0.154367f
C582 variable_delay_unit_4.tristate_inverter_1.en.t0 VSS 0.048564f
C583 variable_delay_unit_4.tristate_inverter_1.en.n1 VSS 0.616703f
C584 variable_delay_unit_4.tristate_inverter_1.en.n2 VSS 0.678061f
C585 variable_delay_unit_4.tristate_inverter_1.en.t7 VSS 0.066961f
C586 variable_delay_unit_4.tristate_inverter_1.en.t3 VSS 0.062029f
C587 variable_delay_unit_4.tristate_inverter_1.en.t5 VSS 0.067187f
C588 variable_delay_unit_4.tristate_inverter_1.en.n3 VSS 0.065756f
C589 variable_delay_unit_4.tristate_inverter_1.en.n4 VSS 0.045654f
C590 variable_delay_unit_1.in.t2 VSS 0.044984f
C591 variable_delay_unit_1.in.t3 VSS 0.017058f
C592 variable_delay_unit_1.in.n0 VSS 0.04731f
C593 variable_delay_unit_1.in.t1 VSS 0.033139f
C594 variable_delay_unit_1.in.t0 VSS 0.105354f
C595 variable_delay_unit_1.in.n1 VSS 0.255341f
C596 variable_delay_unit_1.in.t4 VSS 0.042943f
C597 variable_delay_unit_1.in.t5 VSS 0.013862f
C598 variable_delay_unit_1.in.n2 VSS 0.045159f
C599 variable_delay_unit_1.in.n3 VSS 0.420531f
C600 variable_delay_unit_7.tristate_inverter_1.en.t2 VSS 0.019446f
C601 variable_delay_unit_7.tristate_inverter_1.en.t6 VSS 0.025128f
C602 variable_delay_unit_7.tristate_inverter_1.en.t5 VSS 0.025128f
C603 variable_delay_unit_7.tristate_inverter_1.en.n0 VSS 0.074066f
C604 variable_delay_unit_7.tristate_inverter_1.en.t1 VSS 0.154367f
C605 variable_delay_unit_7.tristate_inverter_1.en.t0 VSS 0.048564f
C606 variable_delay_unit_7.tristate_inverter_1.en.n1 VSS 0.616703f
C607 variable_delay_unit_7.tristate_inverter_1.en.n2 VSS 0.678061f
C608 variable_delay_unit_7.tristate_inverter_1.en.t3 VSS 0.066961f
C609 variable_delay_unit_7.tristate_inverter_1.en.t7 VSS 0.062029f
C610 variable_delay_unit_7.tristate_inverter_1.en.t4 VSS 0.067187f
C611 variable_delay_unit_7.tristate_inverter_1.en.n3 VSS 0.065756f
C612 variable_delay_unit_7.tristate_inverter_1.en.n4 VSS 0.045654f
C613 variable_delay_unit_6.in.t4 VSS 0.044984f
C614 variable_delay_unit_6.in.t5 VSS 0.017058f
C615 variable_delay_unit_6.in.n0 VSS 0.04731f
C616 variable_delay_unit_6.in.t0 VSS 0.033139f
C617 variable_delay_unit_6.in.t1 VSS 0.105354f
C618 variable_delay_unit_6.in.n1 VSS 0.255341f
C619 variable_delay_unit_6.in.t2 VSS 0.042943f
C620 variable_delay_unit_6.in.t3 VSS 0.013862f
C621 variable_delay_unit_6.in.n2 VSS 0.045159f
C622 variable_delay_unit_6.in.n3 VSS 0.420531f
C623 variable_delay_unit_5.in.t4 VSS 0.044984f
C624 variable_delay_unit_5.in.t5 VSS 0.017058f
C625 variable_delay_unit_5.in.n0 VSS 0.04731f
C626 variable_delay_unit_5.in.t0 VSS 0.033139f
C627 variable_delay_unit_5.in.t1 VSS 0.105354f
C628 variable_delay_unit_5.in.n1 VSS 0.255341f
C629 variable_delay_unit_5.in.t2 VSS 0.042943f
C630 variable_delay_unit_5.in.t3 VSS 0.013862f
C631 variable_delay_unit_5.in.n2 VSS 0.045159f
C632 variable_delay_unit_5.in.n3 VSS 0.420531f
C633 variable_delay_unit_0.tristate_inverter_1.en.t4 VSS 0.019446f
C634 variable_delay_unit_0.tristate_inverter_1.en.t2 VSS 0.025128f
C635 variable_delay_unit_0.tristate_inverter_1.en.t6 VSS 0.025128f
C636 variable_delay_unit_0.tristate_inverter_1.en.n0 VSS 0.074066f
C637 variable_delay_unit_0.tristate_inverter_1.en.t1 VSS 0.154367f
C638 variable_delay_unit_0.tristate_inverter_1.en.t0 VSS 0.048564f
C639 variable_delay_unit_0.tristate_inverter_1.en.n1 VSS 0.616703f
C640 variable_delay_unit_0.tristate_inverter_1.en.n2 VSS 0.678061f
C641 variable_delay_unit_0.tristate_inverter_1.en.t5 VSS 0.066961f
C642 variable_delay_unit_0.tristate_inverter_1.en.t7 VSS 0.062029f
C643 variable_delay_unit_0.tristate_inverter_1.en.t3 VSS 0.067187f
C644 variable_delay_unit_0.tristate_inverter_1.en.n3 VSS 0.065756f
C645 variable_delay_unit_0.tristate_inverter_1.en.n4 VSS 0.045654f
C646 variable_delay_unit_1.tristate_inverter_1.en.t5 VSS 0.019446f
C647 variable_delay_unit_1.tristate_inverter_1.en.t2 VSS 0.025128f
C648 variable_delay_unit_1.tristate_inverter_1.en.t3 VSS 0.025128f
C649 variable_delay_unit_1.tristate_inverter_1.en.n0 VSS 0.074066f
C650 variable_delay_unit_1.tristate_inverter_1.en.t1 VSS 0.154367f
C651 variable_delay_unit_1.tristate_inverter_1.en.t0 VSS 0.048564f
C652 variable_delay_unit_1.tristate_inverter_1.en.n1 VSS 0.616703f
C653 variable_delay_unit_1.tristate_inverter_1.en.n2 VSS 0.678061f
C654 variable_delay_unit_1.tristate_inverter_1.en.t7 VSS 0.066961f
C655 variable_delay_unit_1.tristate_inverter_1.en.t4 VSS 0.062029f
C656 variable_delay_unit_1.tristate_inverter_1.en.t6 VSS 0.067187f
C657 variable_delay_unit_1.tristate_inverter_1.en.n3 VSS 0.065756f
C658 variable_delay_unit_1.tristate_inverter_1.en.n4 VSS 0.045654f
C659 variable_delay_unit_2.in.t4 VSS 0.044984f
C660 variable_delay_unit_2.in.t5 VSS 0.017058f
C661 variable_delay_unit_2.in.n0 VSS 0.04731f
C662 variable_delay_unit_2.in.t0 VSS 0.033139f
C663 variable_delay_unit_2.in.t1 VSS 0.105354f
C664 variable_delay_unit_2.in.n1 VSS 0.255341f
C665 variable_delay_unit_2.in.t2 VSS 0.042943f
C666 variable_delay_unit_2.in.t3 VSS 0.013862f
C667 variable_delay_unit_2.in.n2 VSS 0.045159f
C668 variable_delay_unit_2.in.n3 VSS 0.420531f
C669 variable_delay_unit_8.forward.t2 VSS 0.067654f
C670 variable_delay_unit_8.forward.t3 VSS 0.025654f
C671 variable_delay_unit_8.forward.n0 VSS 0.071153f
C672 variable_delay_unit_8.forward.t0 VSS 0.04984f
C673 variable_delay_unit_8.forward.t1 VSS 0.15845f
C674 variable_delay_unit_8.forward.n1 VSS 0.384027f
C675 variable_delay_unit_8.forward.n2 VSS 0.632469f
C676 variable_delay_unit_2.tristate_inverter_1.en.t6 VSS 0.019446f
C677 variable_delay_unit_2.tristate_inverter_1.en.t4 VSS 0.025128f
C678 variable_delay_unit_2.tristate_inverter_1.en.t2 VSS 0.025128f
C679 variable_delay_unit_2.tristate_inverter_1.en.n0 VSS 0.074066f
C680 variable_delay_unit_2.tristate_inverter_1.en.t1 VSS 0.154367f
C681 variable_delay_unit_2.tristate_inverter_1.en.t0 VSS 0.048564f
C682 variable_delay_unit_2.tristate_inverter_1.en.n1 VSS 0.616703f
C683 variable_delay_unit_2.tristate_inverter_1.en.n2 VSS 0.678061f
C684 variable_delay_unit_2.tristate_inverter_1.en.t7 VSS 0.066961f
C685 variable_delay_unit_2.tristate_inverter_1.en.t3 VSS 0.062029f
C686 variable_delay_unit_2.tristate_inverter_1.en.t5 VSS 0.067187f
C687 variable_delay_unit_2.tristate_inverter_1.en.n3 VSS 0.065756f
C688 variable_delay_unit_2.tristate_inverter_1.en.n4 VSS 0.045654f
C689 variable_delay_unit_4.in.t3 VSS 0.044984f
C690 variable_delay_unit_4.in.t5 VSS 0.017058f
C691 variable_delay_unit_4.in.n0 VSS 0.04731f
C692 variable_delay_unit_4.in.t0 VSS 0.033139f
C693 variable_delay_unit_4.in.t1 VSS 0.105354f
C694 variable_delay_unit_4.in.n1 VSS 0.255341f
C695 variable_delay_unit_4.in.t2 VSS 0.042943f
C696 variable_delay_unit_4.in.t4 VSS 0.013862f
C697 variable_delay_unit_4.in.n2 VSS 0.045159f
C698 variable_delay_unit_4.in.n3 VSS 0.420531f
C699 variable_delay_unit_3.in.t4 VSS 0.044984f
C700 variable_delay_unit_3.in.t5 VSS 0.017058f
C701 variable_delay_unit_3.in.n0 VSS 0.04731f
C702 variable_delay_unit_3.in.t1 VSS 0.033139f
C703 variable_delay_unit_3.in.t0 VSS 0.105354f
C704 variable_delay_unit_3.in.n1 VSS 0.255341f
C705 variable_delay_unit_3.in.t2 VSS 0.042943f
C706 variable_delay_unit_3.in.t3 VSS 0.013862f
C707 variable_delay_unit_3.in.n2 VSS 0.045159f
C708 variable_delay_unit_3.in.n3 VSS 0.420531f
C709 variable_delay_unit_8.tristate_inverter_1.en.t4 VSS 0.027086f
C710 variable_delay_unit_8.tristate_inverter_1.en.t2 VSS 0.035f
C711 variable_delay_unit_8.tristate_inverter_1.en.t6 VSS 0.035f
C712 variable_delay_unit_8.tristate_inverter_1.en.n0 VSS 0.103163f
C713 variable_delay_unit_8.tristate_inverter_1.en.t1 VSS 0.215011f
C714 variable_delay_unit_8.tristate_inverter_1.en.t0 VSS 0.067642f
C715 variable_delay_unit_8.tristate_inverter_1.en.n1 VSS 0.85898f
C716 variable_delay_unit_8.tristate_inverter_1.en.n2 VSS 0.944443f
C717 variable_delay_unit_8.tristate_inverter_1.en.t5 VSS 0.093268f
C718 variable_delay_unit_8.tristate_inverter_1.en.t7 VSS 0.086397f
C719 variable_delay_unit_8.tristate_inverter_1.en.t3 VSS 0.093582f
C720 variable_delay_unit_8.tristate_inverter_1.en.n3 VSS 0.091588f
C721 variable_delay_unit_8.tristate_inverter_1.en.n4 VSS 0.06359f
C722 variable_delay_unit_5.tristate_inverter_1.en.t6 VSS 0.019446f
C723 variable_delay_unit_5.tristate_inverter_1.en.t4 VSS 0.025128f
C724 variable_delay_unit_5.tristate_inverter_1.en.t3 VSS 0.025128f
C725 variable_delay_unit_5.tristate_inverter_1.en.n0 VSS 0.074066f
C726 variable_delay_unit_5.tristate_inverter_1.en.t1 VSS 0.154367f
C727 variable_delay_unit_5.tristate_inverter_1.en.t0 VSS 0.048564f
C728 variable_delay_unit_5.tristate_inverter_1.en.n1 VSS 0.616703f
C729 variable_delay_unit_5.tristate_inverter_1.en.n2 VSS 0.678061f
C730 variable_delay_unit_5.tristate_inverter_1.en.t2 VSS 0.066961f
C731 variable_delay_unit_5.tristate_inverter_1.en.t5 VSS 0.062029f
C732 variable_delay_unit_5.tristate_inverter_1.en.t7 VSS 0.067187f
C733 variable_delay_unit_5.tristate_inverter_1.en.n3 VSS 0.065756f
C734 variable_delay_unit_5.tristate_inverter_1.en.n4 VSS 0.045654f
C735 VDD.n0 VSS 0.165217f
C736 VDD.t153 VSS 0.040691f
C737 VDD.n1 VSS 0.042165f
C738 VDD.n2 VSS 0.037662f
C739 VDD.n3 VSS 0.02485f
C740 VDD.t108 VSS 0.169977f
C741 VDD.n4 VSS 0.049067f
C742 VDD.n5 VSS 0.049067f
C743 VDD.t109 VSS 0.040691f
C744 VDD.n6 VSS 0.016963f
C745 VDD.n7 VSS 0.165217f
C746 VDD.n8 VSS 0.046186f
C747 VDD.t33 VSS 0.010843f
C748 VDD.t157 VSS 0.010843f
C749 VDD.n9 VSS 0.031645f
C750 VDD.t49 VSS 0.040033f
C751 VDD.n10 VSS 0.14434f
C752 VDD.n11 VSS 0.062407f
C753 VDD.n12 VSS 0.046186f
C754 VDD.n13 VSS 0.029228f
C755 VDD.n14 VSS 0.159397f
C756 VDD.t114 VSS 0.136186f
C757 VDD.n15 VSS 0.075387f
C758 VDD.n16 VSS 0.075387f
C759 VDD.t85 VSS 0.010843f
C760 VDD.t54 VSS 0.010843f
C761 VDD.n17 VSS 0.031645f
C762 VDD.t58 VSS 0.040033f
C763 VDD.n18 VSS 0.14434f
C764 VDD.t53 VSS 0.077485f
C765 VDD.n19 VSS 0.051657f
C766 VDD.t84 VSS 0.077485f
C767 VDD.t57 VSS 0.152768f
C768 VDD.n20 VSS 0.159397f
C769 VDD.n21 VSS 0.046186f
C770 VDD.n22 VSS 0.165217f
C771 VDD.t161 VSS 0.040691f
C772 VDD.n23 VSS 0.042165f
C773 VDD.n24 VSS 0.037662f
C774 VDD.n25 VSS 0.02485f
C775 VDD.t42 VSS 0.169977f
C776 VDD.n26 VSS 0.049067f
C777 VDD.n27 VSS 0.049067f
C778 VDD.t43 VSS 0.040691f
C779 VDD.n28 VSS 0.016963f
C780 VDD.n29 VSS 0.165217f
C781 VDD.n30 VSS 0.046186f
C782 VDD.t155 VSS 0.010843f
C783 VDD.t102 VSS 0.010843f
C784 VDD.n31 VSS 0.031645f
C785 VDD.t36 VSS 0.040033f
C786 VDD.n32 VSS 0.14434f
C787 VDD.n33 VSS 0.062407f
C788 VDD.n34 VSS 0.046186f
C789 VDD.n35 VSS 0.029228f
C790 VDD.n36 VSS 0.159397f
C791 VDD.t145 VSS 0.136186f
C792 VDD.n37 VSS 0.075387f
C793 VDD.n38 VSS 0.075387f
C794 VDD.t159 VSS 0.010843f
C795 VDD.t139 VSS 0.010843f
C796 VDD.n39 VSS 0.031645f
C797 VDD.t137 VSS 0.040033f
C798 VDD.n40 VSS 0.14434f
C799 VDD.t138 VSS 0.077485f
C800 VDD.n41 VSS 0.051657f
C801 VDD.t158 VSS 0.077485f
C802 VDD.t136 VSS 0.152768f
C803 VDD.n42 VSS 0.159397f
C804 VDD.n43 VSS 0.046186f
C805 VDD.n44 VSS 0.165217f
C806 VDD.t62 VSS 0.040691f
C807 VDD.n45 VSS 0.042165f
C808 VDD.n46 VSS 0.037662f
C809 VDD.n47 VSS 0.02485f
C810 VDD.t142 VSS 0.169977f
C811 VDD.n48 VSS 0.049067f
C812 VDD.n49 VSS 0.049067f
C813 VDD.t143 VSS 0.040691f
C814 VDD.n50 VSS 0.016963f
C815 VDD.n51 VSS 0.165217f
C816 VDD.n52 VSS 0.046186f
C817 VDD.t107 VSS 0.010843f
C818 VDD.t116 VSS 0.010843f
C819 VDD.n53 VSS 0.031645f
C820 VDD.t150 VSS 0.040033f
C821 VDD.n54 VSS 0.14434f
C822 VDD.n55 VSS 0.062407f
C823 VDD.n56 VSS 0.046186f
C824 VDD.n57 VSS 0.029228f
C825 VDD.n58 VSS 0.159397f
C826 VDD.t98 VSS 0.136186f
C827 VDD.n59 VSS 0.075387f
C828 VDD.n60 VSS 0.075387f
C829 VDD.t64 VSS 0.010843f
C830 VDD.t133 VSS 0.010843f
C831 VDD.n61 VSS 0.031645f
C832 VDD.t66 VSS 0.040033f
C833 VDD.n62 VSS 0.14434f
C834 VDD.t132 VSS 0.077485f
C835 VDD.n63 VSS 0.051657f
C836 VDD.t63 VSS 0.077485f
C837 VDD.t65 VSS 0.152768f
C838 VDD.n64 VSS 0.159397f
C839 VDD.n65 VSS 0.046186f
C840 VDD.n66 VSS 0.165217f
C841 VDD.t93 VSS 0.040691f
C842 VDD.n67 VSS 0.042165f
C843 VDD.n68 VSS 0.037662f
C844 VDD.n69 VSS 0.02485f
C845 VDD.t59 VSS 0.169977f
C846 VDD.n70 VSS 0.049067f
C847 VDD.n71 VSS 0.049067f
C848 VDD.t60 VSS 0.040691f
C849 VDD.n72 VSS 0.016963f
C850 VDD.n73 VSS 0.165217f
C851 VDD.n74 VSS 0.046186f
C852 VDD.t97 VSS 0.010843f
C853 VDD.t82 VSS 0.010843f
C854 VDD.n75 VSS 0.031645f
C855 VDD.t41 VSS 0.040033f
C856 VDD.n76 VSS 0.14434f
C857 VDD.n77 VSS 0.062407f
C858 VDD.n78 VSS 0.046186f
C859 VDD.n79 VSS 0.029228f
C860 VDD.n80 VSS 0.159397f
C861 VDD.t6 VSS 0.136186f
C862 VDD.n81 VSS 0.075387f
C863 VDD.n82 VSS 0.075387f
C864 VDD.t47 VSS 0.010843f
C865 VDD.t21 VSS 0.010843f
C866 VDD.n83 VSS 0.031645f
C867 VDD.t19 VSS 0.040033f
C868 VDD.n84 VSS 0.14434f
C869 VDD.t20 VSS 0.077485f
C870 VDD.n85 VSS 0.051657f
C871 VDD.t46 VSS 0.077485f
C872 VDD.t18 VSS 0.152768f
C873 VDD.n86 VSS 0.159397f
C874 VDD.n87 VSS 0.046186f
C875 VDD.n88 VSS 0.165217f
C876 VDD.t1 VSS 0.040691f
C877 VDD.n89 VSS 0.042165f
C878 VDD.n90 VSS 0.037662f
C879 VDD.n91 VSS 0.02485f
C880 VDD.t25 VSS 0.169977f
C881 VDD.n92 VSS 0.049067f
C882 VDD.n93 VSS 0.049067f
C883 VDD.t26 VSS 0.040691f
C884 VDD.n94 VSS 0.016963f
C885 VDD.n95 VSS 0.165217f
C886 VDD.n96 VSS 0.046186f
C887 VDD.t100 VSS 0.010843f
C888 VDD.t52 VSS 0.010843f
C889 VDD.n97 VSS 0.031645f
C890 VDD.t13 VSS 0.040033f
C891 VDD.n98 VSS 0.14434f
C892 VDD.n99 VSS 0.062407f
C893 VDD.n100 VSS 0.046186f
C894 VDD.n101 VSS 0.029228f
C895 VDD.n102 VSS 0.159397f
C896 VDD.t37 VSS 0.136186f
C897 VDD.n103 VSS 0.075387f
C898 VDD.n104 VSS 0.075387f
C899 VDD.t3 VSS 0.010843f
C900 VDD.t56 VSS 0.010843f
C901 VDD.n105 VSS 0.031645f
C902 VDD.t68 VSS 0.040033f
C903 VDD.n106 VSS 0.14434f
C904 VDD.t55 VSS 0.077485f
C905 VDD.n107 VSS 0.051657f
C906 VDD.t2 VSS 0.077485f
C907 VDD.t67 VSS 0.152768f
C908 VDD.n108 VSS 0.159397f
C909 VDD.n109 VSS 0.046186f
C910 VDD.n110 VSS 0.165217f
C911 VDD.t141 VSS 0.040691f
C912 VDD.n111 VSS 0.042165f
C913 VDD.n112 VSS 0.037662f
C914 VDD.n113 VSS 0.02485f
C915 VDD.t30 VSS 0.169977f
C916 VDD.n114 VSS 0.049067f
C917 VDD.n115 VSS 0.049067f
C918 VDD.t31 VSS 0.040691f
C919 VDD.n116 VSS 0.016963f
C920 VDD.n117 VSS 0.165217f
C921 VDD.n118 VSS 0.046186f
C922 VDD.t118 VSS 0.010843f
C923 VDD.t135 VSS 0.010843f
C924 VDD.n119 VSS 0.031645f
C925 VDD.t23 VSS 0.040033f
C926 VDD.n120 VSS 0.14434f
C927 VDD.n121 VSS 0.062407f
C928 VDD.n122 VSS 0.046186f
C929 VDD.n123 VSS 0.029228f
C930 VDD.n124 VSS 0.159397f
C931 VDD.t105 VSS 0.136186f
C932 VDD.n125 VSS 0.075387f
C933 VDD.n126 VSS 0.075387f
C934 VDD.t28 VSS 0.010843f
C935 VDD.t17 VSS 0.010843f
C936 VDD.n127 VSS 0.031645f
C937 VDD.t91 VSS 0.040033f
C938 VDD.n128 VSS 0.14434f
C939 VDD.t16 VSS 0.077485f
C940 VDD.n129 VSS 0.051657f
C941 VDD.t27 VSS 0.077485f
C942 VDD.t90 VSS 0.152768f
C943 VDD.n130 VSS 0.159397f
C944 VDD.n131 VSS 0.046186f
C945 VDD.n132 VSS 0.165217f
C946 VDD.t39 VSS 0.040691f
C947 VDD.n133 VSS 0.042165f
C948 VDD.n134 VSS 0.037662f
C949 VDD.n135 VSS 0.02485f
C950 VDD.t86 VSS 0.169977f
C951 VDD.n136 VSS 0.049067f
C952 VDD.n137 VSS 0.049067f
C953 VDD.t87 VSS 0.040691f
C954 VDD.n138 VSS 0.016963f
C955 VDD.n139 VSS 0.165217f
C956 VDD.n140 VSS 0.046186f
C957 VDD.t95 VSS 0.010843f
C958 VDD.t148 VSS 0.010843f
C959 VDD.n141 VSS 0.031645f
C960 VDD.t124 VSS 0.040033f
C961 VDD.n142 VSS 0.14434f
C962 VDD.n143 VSS 0.062407f
C963 VDD.n144 VSS 0.046186f
C964 VDD.n145 VSS 0.029228f
C965 VDD.n146 VSS 0.159397f
C966 VDD.t50 VSS 0.136186f
C967 VDD.n147 VSS 0.075387f
C968 VDD.n148 VSS 0.075387f
C969 VDD.t113 VSS 0.010843f
C970 VDD.t128 VSS 0.010843f
C971 VDD.n149 VSS 0.031645f
C972 VDD.t126 VSS 0.040033f
C973 VDD.n150 VSS 0.14434f
C974 VDD.t127 VSS 0.077485f
C975 VDD.n151 VSS 0.051657f
C976 VDD.t112 VSS 0.077485f
C977 VDD.t125 VSS 0.152768f
C978 VDD.n152 VSS 0.159397f
C979 VDD.n153 VSS 0.046186f
C980 VDD.n154 VSS 0.165217f
C981 VDD.t80 VSS 0.040691f
C982 VDD.n155 VSS 0.042165f
C983 VDD.n156 VSS 0.037662f
C984 VDD.n157 VSS 0.02485f
C985 VDD.t162 VSS 0.169977f
C986 VDD.n158 VSS 0.049067f
C987 VDD.n159 VSS 0.049067f
C988 VDD.t163 VSS 0.040691f
C989 VDD.n160 VSS 0.016963f
C990 VDD.n161 VSS 0.165217f
C991 VDD.n162 VSS 0.046186f
C992 VDD.t11 VSS 0.010843f
C993 VDD.t15 VSS 0.010843f
C994 VDD.n163 VSS 0.031645f
C995 VDD.t122 VSS 0.040033f
C996 VDD.n164 VSS 0.14434f
C997 VDD.n165 VSS 0.062407f
C998 VDD.n166 VSS 0.046186f
C999 VDD.n167 VSS 0.029228f
C1000 VDD.n168 VSS 0.159397f
C1001 VDD.t34 VSS 0.136186f
C1002 VDD.n169 VSS 0.075387f
C1003 VDD.n170 VSS 0.075387f
C1004 VDD.t77 VSS 0.010843f
C1005 VDD.t74 VSS 0.010843f
C1006 VDD.n171 VSS 0.031645f
C1007 VDD.t71 VSS 0.040033f
C1008 VDD.n172 VSS 0.14434f
C1009 VDD.t73 VSS 0.077485f
C1010 VDD.n173 VSS 0.051657f
C1011 VDD.t76 VSS 0.077485f
C1012 VDD.t70 VSS 0.152768f
C1013 VDD.n174 VSS 0.159397f
C1014 VDD.n175 VSS 0.046294f
C1015 VDD.n176 VSS 0.029054f
C1016 VDD.n177 VSS 0.02704f
C1017 VDD.n178 VSS 0.062407f
C1018 VDD.n179 VSS 0.046186f
C1019 VDD.n180 VSS 0.029228f
C1020 VDD.n181 VSS 0.278242f
C1021 VDD.n182 VSS 0.278242f
C1022 VDD.t129 VSS 0.136186f
C1023 VDD.t10 VSS 0.077485f
C1024 VDD.t121 VSS 0.152768f
C1025 VDD.t14 VSS 0.077485f
C1026 VDD.n183 VSS 0.051657f
C1027 VDD.n184 VSS 0.075387f
C1028 VDD.n185 VSS 0.075387f
C1029 VDD.n186 VSS 0.02704f
C1030 VDD.n187 VSS 0.029353f
C1031 VDD.n188 VSS 0.035307f
C1032 VDD.n189 VSS 0.058679f
C1033 VDD.n190 VSS 0.011306f
C1034 VDD.n191 VSS 0.075071f
C1035 VDD.n192 VSS 0.039533f
C1036 VDD.n193 VSS 0.037662f
C1037 VDD.n194 VSS 0.02485f
C1038 VDD.n195 VSS 0.134954f
C1039 VDD.n196 VSS 0.134954f
C1040 VDD.t79 VSS 0.169977f
C1041 VDD.n197 VSS 0.016963f
C1042 VDD.n198 VSS 0.049067f
C1043 VDD.n199 VSS 0.049067f
C1044 VDD.n200 VSS 0.011306f
C1045 VDD.n201 VSS 0.075071f
C1046 VDD.n202 VSS 0.041088f
C1047 VDD.t169 VSS 0.005122f
C1048 VDD.t168 VSS 0.006619f
C1049 VDD.t166 VSS 0.006619f
C1050 VDD.n203 VSS 0.01951f
C1051 VDD.t75 VSS 0.016339f
C1052 VDD.t69 VSS 0.017698f
C1053 VDD.n204 VSS 0.017321f
C1054 VDD.t72 VSS 0.017638f
C1055 VDD.n205 VSS 0.012026f
C1056 VDD.n206 VSS 0.126355f
C1057 VDD.n207 VSS 0.100414f
C1058 VDD.t78 VSS 0.016563f
C1059 VDD.t167 VSS 0.005347f
C1060 VDD.n208 VSS 0.016305f
C1061 VDD.n209 VSS 0.11626f
C1062 VDD.n210 VSS 0.037036f
C1063 VDD.n211 VSS 0.029624f
C1064 VDD.n212 VSS 0.029054f
C1065 VDD.n213 VSS 0.02704f
C1066 VDD.n214 VSS 0.062407f
C1067 VDD.n215 VSS 0.046186f
C1068 VDD.n216 VSS 0.029228f
C1069 VDD.n217 VSS 0.278242f
C1070 VDD.n218 VSS 0.278242f
C1071 VDD.t165 VSS 0.136186f
C1072 VDD.t94 VSS 0.077485f
C1073 VDD.t123 VSS 0.152768f
C1074 VDD.t147 VSS 0.077485f
C1075 VDD.n219 VSS 0.051657f
C1076 VDD.n220 VSS 0.075387f
C1077 VDD.n221 VSS 0.075387f
C1078 VDD.n222 VSS 0.02704f
C1079 VDD.n223 VSS 0.029353f
C1080 VDD.n224 VSS 0.035307f
C1081 VDD.n225 VSS 0.058679f
C1082 VDD.n226 VSS 0.011306f
C1083 VDD.n227 VSS 0.075071f
C1084 VDD.n228 VSS 0.039533f
C1085 VDD.n229 VSS 0.037662f
C1086 VDD.n230 VSS 0.02485f
C1087 VDD.n231 VSS 0.134954f
C1088 VDD.n232 VSS 0.134954f
C1089 VDD.t38 VSS 0.169977f
C1090 VDD.n233 VSS 0.016963f
C1091 VDD.n234 VSS 0.049067f
C1092 VDD.n235 VSS 0.049067f
C1093 VDD.n236 VSS 0.011306f
C1094 VDD.n237 VSS 0.075071f
C1095 VDD.n238 VSS 0.066742f
C1096 VDD.n239 VSS 0.029624f
C1097 VDD.n240 VSS 0.029054f
C1098 VDD.n241 VSS 0.02704f
C1099 VDD.n242 VSS 0.062407f
C1100 VDD.n243 VSS 0.046186f
C1101 VDD.n244 VSS 0.029228f
C1102 VDD.n245 VSS 0.278242f
C1103 VDD.n246 VSS 0.278242f
C1104 VDD.t164 VSS 0.136186f
C1105 VDD.t117 VSS 0.077485f
C1106 VDD.t22 VSS 0.152768f
C1107 VDD.t134 VSS 0.077485f
C1108 VDD.n247 VSS 0.051657f
C1109 VDD.n248 VSS 0.075387f
C1110 VDD.n249 VSS 0.075387f
C1111 VDD.n250 VSS 0.02704f
C1112 VDD.n251 VSS 0.029353f
C1113 VDD.n252 VSS 0.035307f
C1114 VDD.n253 VSS 0.058679f
C1115 VDD.n254 VSS 0.011306f
C1116 VDD.n255 VSS 0.075071f
C1117 VDD.n256 VSS 0.039533f
C1118 VDD.n257 VSS 0.037662f
C1119 VDD.n258 VSS 0.02485f
C1120 VDD.n259 VSS 0.134954f
C1121 VDD.n260 VSS 0.134954f
C1122 VDD.t140 VSS 0.169977f
C1123 VDD.n261 VSS 0.016963f
C1124 VDD.n262 VSS 0.049067f
C1125 VDD.n263 VSS 0.049067f
C1126 VDD.n264 VSS 0.011306f
C1127 VDD.n265 VSS 0.075071f
C1128 VDD.n266 VSS 0.066742f
C1129 VDD.n267 VSS 0.029624f
C1130 VDD.n268 VSS 0.029054f
C1131 VDD.n269 VSS 0.02704f
C1132 VDD.n270 VSS 0.062407f
C1133 VDD.n271 VSS 0.046186f
C1134 VDD.n272 VSS 0.029228f
C1135 VDD.n273 VSS 0.278242f
C1136 VDD.n274 VSS 0.278242f
C1137 VDD.t29 VSS 0.136186f
C1138 VDD.t99 VSS 0.077485f
C1139 VDD.t12 VSS 0.152768f
C1140 VDD.t51 VSS 0.077485f
C1141 VDD.n275 VSS 0.051657f
C1142 VDD.n276 VSS 0.075387f
C1143 VDD.n277 VSS 0.075387f
C1144 VDD.n278 VSS 0.02704f
C1145 VDD.n279 VSS 0.029353f
C1146 VDD.n280 VSS 0.035307f
C1147 VDD.n281 VSS 0.058679f
C1148 VDD.n282 VSS 0.011306f
C1149 VDD.n283 VSS 0.075071f
C1150 VDD.n284 VSS 0.039533f
C1151 VDD.n285 VSS 0.037662f
C1152 VDD.n286 VSS 0.02485f
C1153 VDD.n287 VSS 0.134954f
C1154 VDD.n288 VSS 0.134954f
C1155 VDD.t0 VSS 0.169977f
C1156 VDD.n289 VSS 0.016963f
C1157 VDD.n290 VSS 0.049067f
C1158 VDD.n291 VSS 0.049067f
C1159 VDD.n292 VSS 0.011306f
C1160 VDD.n293 VSS 0.075071f
C1161 VDD.n294 VSS 0.066742f
C1162 VDD.n295 VSS 0.029624f
C1163 VDD.n296 VSS 0.029054f
C1164 VDD.n297 VSS 0.02704f
C1165 VDD.n298 VSS 0.062407f
C1166 VDD.n299 VSS 0.046186f
C1167 VDD.n300 VSS 0.029228f
C1168 VDD.n301 VSS 0.278242f
C1169 VDD.n302 VSS 0.278242f
C1170 VDD.t24 VSS 0.136186f
C1171 VDD.t96 VSS 0.077485f
C1172 VDD.t40 VSS 0.152768f
C1173 VDD.t81 VSS 0.077485f
C1174 VDD.n303 VSS 0.051657f
C1175 VDD.n304 VSS 0.075387f
C1176 VDD.n305 VSS 0.075387f
C1177 VDD.n306 VSS 0.02704f
C1178 VDD.n307 VSS 0.029353f
C1179 VDD.n308 VSS 0.035307f
C1180 VDD.n309 VSS 0.058679f
C1181 VDD.n310 VSS 0.011306f
C1182 VDD.n311 VSS 0.075071f
C1183 VDD.n312 VSS 0.039533f
C1184 VDD.n313 VSS 0.037662f
C1185 VDD.n314 VSS 0.02485f
C1186 VDD.n315 VSS 0.134954f
C1187 VDD.n316 VSS 0.134954f
C1188 VDD.t92 VSS 0.169977f
C1189 VDD.n317 VSS 0.016963f
C1190 VDD.n318 VSS 0.049067f
C1191 VDD.n319 VSS 0.049067f
C1192 VDD.n320 VSS 0.011306f
C1193 VDD.n321 VSS 0.075071f
C1194 VDD.n322 VSS 0.066742f
C1195 VDD.n323 VSS 0.029624f
C1196 VDD.n324 VSS 0.029054f
C1197 VDD.n325 VSS 0.02704f
C1198 VDD.n326 VSS 0.062407f
C1199 VDD.n327 VSS 0.046186f
C1200 VDD.n328 VSS 0.029228f
C1201 VDD.n329 VSS 0.278242f
C1202 VDD.n330 VSS 0.278242f
C1203 VDD.t144 VSS 0.136186f
C1204 VDD.t106 VSS 0.077485f
C1205 VDD.t149 VSS 0.152768f
C1206 VDD.t115 VSS 0.077485f
C1207 VDD.n331 VSS 0.051657f
C1208 VDD.n332 VSS 0.075387f
C1209 VDD.n333 VSS 0.075387f
C1210 VDD.n334 VSS 0.02704f
C1211 VDD.n335 VSS 0.029353f
C1212 VDD.n336 VSS 0.035307f
C1213 VDD.n337 VSS 0.058679f
C1214 VDD.n338 VSS 0.011306f
C1215 VDD.n339 VSS 0.075071f
C1216 VDD.n340 VSS 0.039533f
C1217 VDD.n341 VSS 0.037662f
C1218 VDD.n342 VSS 0.02485f
C1219 VDD.n343 VSS 0.134954f
C1220 VDD.n344 VSS 0.134954f
C1221 VDD.t61 VSS 0.169977f
C1222 VDD.n345 VSS 0.016963f
C1223 VDD.n346 VSS 0.049067f
C1224 VDD.n347 VSS 0.049067f
C1225 VDD.n348 VSS 0.011306f
C1226 VDD.n349 VSS 0.075071f
C1227 VDD.n350 VSS 0.066742f
C1228 VDD.n351 VSS 0.029624f
C1229 VDD.n352 VSS 0.029054f
C1230 VDD.n353 VSS 0.02704f
C1231 VDD.n354 VSS 0.062407f
C1232 VDD.n355 VSS 0.046186f
C1233 VDD.n356 VSS 0.029228f
C1234 VDD.n357 VSS 0.278242f
C1235 VDD.n358 VSS 0.278242f
C1236 VDD.t83 VSS 0.136186f
C1237 VDD.t154 VSS 0.077485f
C1238 VDD.t35 VSS 0.152768f
C1239 VDD.t101 VSS 0.077485f
C1240 VDD.n359 VSS 0.051657f
C1241 VDD.n360 VSS 0.075387f
C1242 VDD.n361 VSS 0.075387f
C1243 VDD.n362 VSS 0.02704f
C1244 VDD.n363 VSS 0.029353f
C1245 VDD.n364 VSS 0.035307f
C1246 VDD.n365 VSS 0.058679f
C1247 VDD.n366 VSS 0.011306f
C1248 VDD.n367 VSS 0.075071f
C1249 VDD.n368 VSS 0.039533f
C1250 VDD.n369 VSS 0.037662f
C1251 VDD.n370 VSS 0.02485f
C1252 VDD.n371 VSS 0.134954f
C1253 VDD.n372 VSS 0.134954f
C1254 VDD.t160 VSS 0.169977f
C1255 VDD.n373 VSS 0.016963f
C1256 VDD.n374 VSS 0.049067f
C1257 VDD.n375 VSS 0.049067f
C1258 VDD.n376 VSS 0.011306f
C1259 VDD.n377 VSS 0.075071f
C1260 VDD.n378 VSS 0.066742f
C1261 VDD.n379 VSS 0.029624f
C1262 VDD.n380 VSS 0.029054f
C1263 VDD.n381 VSS 0.02704f
C1264 VDD.n382 VSS 0.062407f
C1265 VDD.n383 VSS 0.046186f
C1266 VDD.n384 VSS 0.029228f
C1267 VDD.n385 VSS 0.278242f
C1268 VDD.n386 VSS 0.278242f
C1269 VDD.t146 VSS 0.136186f
C1270 VDD.t32 VSS 0.077485f
C1271 VDD.t48 VSS 0.152768f
C1272 VDD.t156 VSS 0.077485f
C1273 VDD.n387 VSS 0.051657f
C1274 VDD.n388 VSS 0.075387f
C1275 VDD.n389 VSS 0.075387f
C1276 VDD.n390 VSS 0.02704f
C1277 VDD.n391 VSS 0.029353f
C1278 VDD.n392 VSS 0.035307f
C1279 VDD.n393 VSS 0.058679f
C1280 VDD.n394 VSS 0.011306f
C1281 VDD.n395 VSS 0.075071f
C1282 VDD.n396 VSS 0.039533f
C1283 VDD.n397 VSS 0.037662f
C1284 VDD.n398 VSS 0.02485f
C1285 VDD.n399 VSS 0.134954f
C1286 VDD.n400 VSS 0.134954f
C1287 VDD.t152 VSS 0.169977f
C1288 VDD.n401 VSS 0.016963f
C1289 VDD.n402 VSS 0.049067f
C1290 VDD.n403 VSS 0.049067f
C1291 VDD.n404 VSS 0.011306f
C1292 VDD.n405 VSS 0.075071f
C1293 VDD.n406 VSS 0.066742f
C1294 VDD.n407 VSS 0.046186f
C1295 VDD.t111 VSS 0.010843f
C1296 VDD.t8 VSS 0.010843f
C1297 VDD.n408 VSS 0.031645f
C1298 VDD.t131 VSS 0.040033f
C1299 VDD.n409 VSS 0.14434f
C1300 VDD.n410 VSS 0.062407f
C1301 VDD.n411 VSS 0.075387f
C1302 VDD.n412 VSS 0.159397f
C1303 VDD.t130 VSS 0.152768f
C1304 VDD.t110 VSS 0.077485f
C1305 VDD.n413 VSS 0.051657f
C1306 VDD.t7 VSS 0.077485f
C1307 VDD.t151 VSS 0.136186f
C1308 VDD.t9 VSS 0.136186f
C1309 VDD.n414 VSS 0.075387f
C1310 VDD.n415 VSS 0.075387f
C1311 VDD.t104 VSS 0.010843f
C1312 VDD.t120 VSS 0.010843f
C1313 VDD.n416 VSS 0.031645f
C1314 VDD.t45 VSS 0.040033f
C1315 VDD.n417 VSS 0.14434f
C1316 VDD.t103 VSS 0.077485f
C1317 VDD.n418 VSS 0.051657f
C1318 VDD.t119 VSS 0.077485f
C1319 VDD.t44 VSS 0.152768f
C1320 VDD.n419 VSS 0.159397f
C1321 VDD.n420 VSS 0.046186f
C1322 VDD.n421 VSS 0.165217f
C1323 VDD.t5 VSS 0.040691f
C1324 VDD.n422 VSS 0.075071f
C1325 VDD.n423 VSS 0.049067f
C1326 VDD.n424 VSS 0.02485f
C1327 VDD.n425 VSS 0.037662f
C1328 VDD.t89 VSS 0.040691f
C1329 VDD.n426 VSS 0.075071f
C1330 VDD.n427 VSS 0.049067f
C1331 VDD.n428 VSS 0.062674f
C1332 VDD.n429 VSS 0.016963f
C1333 VDD.t4 VSS 0.169977f
C1334 VDD.n430 VSS 0.134954f
C1335 VDD.n431 VSS 0.02485f
C1336 VDD.n432 VSS 0.134954f
C1337 VDD.t88 VSS 0.169977f
C1338 VDD.n433 VSS 0.016963f
C1339 VDD.n434 VSS 0.165217f
C1340 VDD.n435 VSS 0.049067f
C1341 VDD.n436 VSS 0.011306f
C1342 VDD.n437 VSS 0.042165f
C1343 VDD.n438 VSS 0.039533f
C1344 VDD.n439 VSS 0.037662f
C1345 VDD.n440 VSS 0.049067f
C1346 VDD.n441 VSS 0.011306f
C1347 VDD.n442 VSS 0.058679f
C1348 VDD.n443 VSS 0.035307f
C1349 VDD.n444 VSS 0.029353f
C1350 VDD.n445 VSS 0.02704f
C1351 VDD.n446 VSS 0.062407f
C1352 VDD.n447 VSS 0.046186f
C1353 VDD.n448 VSS 0.029228f
C1354 VDD.n449 VSS 0.278242f
C1355 VDD.n450 VSS 0.278242f
C1356 VDD.n451 VSS 0.029228f
C1357 VDD.n452 VSS 0.046186f
C1358 VDD.n453 VSS 0.075387f
C1359 VDD.n454 VSS 0.02704f
C1360 VDD.n455 VSS 0.029054f
C1361 VDD.n456 VSS 0.029624f
.ends

