* NGSPICE file created from fine_delay_unit_parax.ext - technology: sky130A

.subckt fine_delay_unit_parax in t0 t1 out VDD VSS
X0 a_544_434# in.t0 a_632_434# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X1 a_896_n120# in.t1 a_632_434# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X2 a_544_434# in.t2 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X3 VSS.t8 t1.t0 a_896_n120# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X4 out.t0 a_544_434# VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X5 a_632_434# in.t3 a_544_434# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X6 a_632_434# in.t4 a_544_434# VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X7 VSS.t3 in.t5 a_896_n120# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X8 out.t1 a_544_434# VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X9 a_896_n120# t0.t0 a_632_434# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
R0 in in.t2 757.207
R1 in.n2 in.t4 343.827
R2 in.n0 in.t5 343.827
R3 in.n2 in.t0 202.44
R4 in.n0 in.t1 202.44
R5 in.n1 in.t3 202.44
R6 in in.n3 167.328
R7 in.n1 in.n0 141.387
R8 in.n3 in.n2 41.7738
R9 in.n3 in.n1 41.7738
R10 VSS.n11 VSS.n8 4447.27
R11 VSS.n14 VSS.n11 3442.57
R12 VSS.n8 VSS.n5 3165.68
R13 VSS.n17 VSS.n7 1438.1
R14 VSS.n17 VSS.n5 1065.44
R15 VSS.t0 VSS.n8 559.691
R16 VSS.n15 VSS.n14 348.32
R17 VSS.t2 VSS.t0 303.449
R18 VSS.t6 VSS.t2 303.449
R19 VSS.t5 VSS.t7 303.449
R20 VSS.n7 VSS.n6 292.5
R21 VSS.n12 VSS.n4 288.961
R22 VSS.n16 VSS.t4 286.207
R23 VSS.n13 VSS.n12 223.68
R24 VSS.n15 VSS.n7 217.493
R25 VSS.n19 VSS.n4 205.69
R26 VSS.n10 VSS.t6 155.173
R27 VSS.t4 VSS.n15 149.625
R28 VSS.n18 VSS.n17 146.25
R29 VSS.n17 VSS.n16 146.25
R30 VSS.n13 VSS.n6 143.361
R31 VSS.n18 VSS.n6 93.4405
R32 VSS.n9 VSS.t5 93.1039
R33 VSS.n19 VSS.n18 69.2272
R34 VSS.n2 VSS.n1 67.5509
R35 VSS.n12 VSS.n11 65.0005
R36 VSS.n11 VSS.n10 65.0005
R37 VSS.n14 VSS.n13 65.0005
R38 VSS.n10 VSS.n9 55.1729
R39 VSS.n2 VSS.t8 41.3938
R40 VSS.n8 VSS.n4 39.0005
R41 VSS.n19 VSS.n5 24.3755
R42 VSS.n9 VSS.n5 24.3755
R43 VSS.n1 VSS.t1 17.4005
R44 VSS.n1 VSS.t3 17.4005
R45 VSS.n16 VSS.t7 17.2419
R46 VSS.n13 VSS.n0 2.913
R47 VSS.n18 VSS.n0 2.3255
R48 VSS.n4 VSS.n3 2.12011
R49 VSS.n3 VSS.n2 0.957022
R50 VSS.n21 VSS.n0 0.440404
R51 VSS.n20 VSS.n19 0.423227
R52 VSS VSS.n21 0.306056
R53 VSS.n20 VSS.n3 0.168035
R54 VSS.n21 VSS.n20 0.104667
R55 VDD.n6 VDD.n3 1271.17
R56 VDD.n8 VDD.n3 408.981
R57 VDD.n11 VDD.n10 313.632
R58 VDD.n5 VDD.n2 135.591
R59 VDD.n12 VDD.n0 129.013
R60 VDD.n4 VDD.t1 84.7771
R61 VDD.n14 VDD.t3 84.7716
R62 VDD.n11 VDD.n3 61.6672
R63 VDD.n7 VDD.n2 43.625
R64 VDD.n10 VDD.n0 35.5275
R65 VDD.n9 VDD.t2 20.8338
R66 VDD.n8 VDD.n7 20.5561
R67 VDD.n9 VDD.n8 20.5561
R68 VDD.n6 VDD.n5 20.5561
R69 VDD.n9 VDD.n6 20.5561
R70 VDD.n12 VDD.n11 7.70883
R71 VDD.n12 VDD.n2 6.57828
R72 VDD.n10 VDD.n9 5.33119
R73 VDD.n5 VDD.n4 2.13168
R74 VDD.t2 VDD.t0 2.08383
R75 VDD.n15 VDD.n0 1.96588
R76 VDD.n7 VDD.n1 1.54255
R77 VDD.n13 VDD.n12 0.423227
R78 VDD VDD.n15 0.182792
R79 VDD.n14 VDD.n13 0.127236
R80 VDD.n4 VDD.n1 0.115083
R81 VDD.n15 VDD.n14 0.0899097
R82 VDD.n13 VDD.n1 0.0647361
R83 t1 t1.t0 727.149
R84 out out.t1 84.8857
R85 out out.t0 84.6628
R86 t0 t0.t0 577.703
C0 a_896_n120# out 7.3e-20
C1 t1 out 0.034216f
C2 in a_632_434# 0.244525f
C3 VDD t1 0.004852f
C4 t0 in 0.009158f
C5 t0 a_632_434# 0.022005f
C6 a_544_434# out 0.115353f
C7 VDD a_544_434# 1.2503f
C8 a_896_n120# t1 0.013742f
C9 out in 0.002069f
C10 out a_632_434# 3.44e-20
C11 a_544_434# a_896_n120# 0.019821f
C12 a_544_434# t1 0.010812f
C13 VDD in 0.275771f
C14 t0 VDD 4.29e-19
C15 a_896_n120# in 0.028846f
C16 a_896_n120# a_632_434# 0.556904f
C17 t1 in 0.020481f
C18 t1 a_632_434# 0.001628f
C19 t0 a_896_n120# 0.02185f
C20 t0 t1 0.014805f
C21 VDD out 0.963042f
C22 a_544_434# in 0.250047f
C23 a_544_434# a_632_434# 0.53267f
C24 t0 a_544_434# 0.003337f
C25 t0 VSS 0.314637f
C26 t1 VSS 0.377692f
C27 out VSS 0.493979f
C28 in VSS 1.07559f
C29 VDD VSS 3.80486f
C30 a_896_n120# VSS 0.612975f
C31 a_632_434# VSS 0.387205f
C32 a_544_434# VSS 0.745736f
.ends

