magic
tech sky130A
timestamp 1731213143
<< end >>
