* NGSPICE file created from input_stage.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_6H9P4D a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
**devattr s=11600,516 d=11600,516
.ends

.subckt sky130_fd_pr__pfet_01v8_2K9SAN a_n73_n300# w_n109_n362# a_15_n300# a_n15_n326#
X0 a_15_n300# a_n15_n326# a_n73_n300# w_n109_n362# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
**devattr s=34800,1316 d=34800,1316
.ends

.subckt sky130_fd_pr__nfet_01v8_TC9PQS a_15_n200# a_n15_n226# a_n73_n200# VSUBS
X0 a_15_n200# a_n15_n226# a_n73_n200# VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
**devattr s=23200,916 d=23200,916
.ends

.subckt fine_delay_unit in t0 t1 out VDD VSS
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 a_978_702# m1_814_280# in VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_1 m1_814_280# a_978_702# in VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__pfet_01v8_2K9SAN_0 VDD VDD a_978_702# in sky130_fd_pr__pfet_01v8_2K9SAN
Xsky130_fd_pr__nfet_01v8_6H9P4D_2 a_978_702# m1_814_280# in VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__pfet_01v8_2K9SAN_1 VDD VDD out a_978_702# sky130_fd_pr__pfet_01v8_2K9SAN
Xsky130_fd_pr__nfet_01v8_6H9P4D_3 m1_814_280# m1_902_280# in VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_4 m1_902_280# VSS in VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_6H9P4D_5 VSS out a_978_702# VSS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__nfet_01v8_TC9PQS_0 m1_902_280# t0 m1_814_280# VSS sky130_fd_pr__nfet_01v8_TC9PQS
Xsky130_fd_pr__nfet_01v8_TC9PQS_1 VSS t1 m1_902_280# VSS sky130_fd_pr__nfet_01v8_TC9PQS
.ends

.subckt inverter_3_1 w_30_230# m1_250_162# sky130_fd_pr__pfet_01v8_2K9SAN_0/VSUBS
+ a_136_200#
Xsky130_fd_pr__nfet_01v8_6H9P4D_0 sky130_fd_pr__pfet_01v8_2K9SAN_0/VSUBS m1_250_162#
+ a_136_200# sky130_fd_pr__pfet_01v8_2K9SAN_0/VSUBS sky130_fd_pr__nfet_01v8_6H9P4D
Xsky130_fd_pr__pfet_01v8_2K9SAN_0 w_30_230# w_30_230# m1_250_162# a_136_200# sky130_fd_pr__pfet_01v8_2K9SAN
.ends

.subckt nand_gate a b out VDD VSS
Xsky130_fd_pr__pfet_01v8_2K9SAN_0 VDD VDD out a sky130_fd_pr__pfet_01v8_2K9SAN
Xsky130_fd_pr__pfet_01v8_2K9SAN_1 out VDD VDD b sky130_fd_pr__pfet_01v8_2K9SAN
Xsky130_fd_pr__nfet_01v8_TC9PQS_0 sky130_fd_pr__nfet_01v8_TC9PQS_0/a_15_n200# a out
+ VSS sky130_fd_pr__nfet_01v8_TC9PQS
Xsky130_fd_pr__nfet_01v8_TC9PQS_1 VSS b sky130_fd_pr__nfet_01v8_TC9PQS_0/a_15_n200#
+ VSS sky130_fd_pr__nfet_01v8_TC9PQS
.ends

.subckt input_stage in en t0 t1 t2 t3 out VDD VSS
Xfine_delay_unit_0 fine_delay_unit_0/in t0 t1 fine_delay_unit_1/in VDD VSS fine_delay_unit
Xfine_delay_unit_1 fine_delay_unit_1/in t2 t3 out VDD VSS fine_delay_unit
Xinverter_3_1_0 VDD fine_delay_unit_0/in VSS nand_gate_0/out inverter_3_1
Xnand_gate_0 en in nand_gate_0/out VDD VSS nand_gate
.ends

