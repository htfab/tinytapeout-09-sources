* NGSPICE file created from variable_delay_short_parax.ext - technology: sky130A

.subckt variable_delay_short_parax in en_1 out en_2 en_3 en_0 en_4 VSS VDD
X0 a_16354_772# variable_delay_unit_5.tristate_inverter_1.en.t2 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X1 VDD.t54 en_1.t0 a_5444_772# VDD.t53 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X2 VSS.t71 variable_delay_unit_2.tristate_inverter_1.en.t2 a_8392_352# VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X3 variable_delay_unit_4.in.t1 variable_delay_unit_3.in.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X4 a_16354_352# VDD.t112 VSS.t79 VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X5 VDD.t24 en_1.t1 a_5444_772# VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X6 variable_delay_unit_3.in.t1 variable_delay_unit_2.in.t2 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X7 VDD.t50 en_0.t0 a_2496_772# VDD.t49 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X8 VDD.t80 VDD.t78 a_17236_772# VDD.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X9 variable_delay_unit_4.in.t0 variable_delay_unit_3.in.t3 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X10 VSS.t36 variable_delay_unit_1.tristate_inverter_1.en.t2 a_5444_352# VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X11 variable_delay_unit_3.in.t0 variable_delay_unit_2.in.t3 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 VSS.t48 variable_delay_unit_1.tristate_inverter_1.en.t3 a_5444_352# VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X13 VSS.t85 variable_delay_unit_5.tristate_inverter_1.en.t3 a_17236_352# VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X14 VDD.t94 variable_delay_unit_2.tristate_inverter_1.en.t3 a_7510_772# VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X15 VSS.t50 variable_delay_unit_0.tristate_inverter_1.en.t2 a_2496_352# VSS.t49 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X16 variable_delay_unit_1.out variable_delay_unit_2.in.t4 a_4562_772# VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X17 variable_delay_unit_5.forward.t1 variable_delay_unit_5.in.t2 VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X18 VDD.t57 en_4.t0 a_14288_772# VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X19 VDD.t108 variable_delay_unit_1.tristate_inverter_1.en.t4 a_4562_772# VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X20 VDD.t52 en_3.t0 a_11340_772# VDD.t51 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X21 variable_delay_unit_0.tristate_inverter_1.en.t1 en_0.t1 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X22 VSS.t7 en_2.t0 a_7510_352# VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X23 variable_delay_unit_1.out variable_delay_unit_2.in.t5 a_4562_352# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X24 out.t2 variable_delay_unit_1.in.t2 a_1614_772# VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X25 variable_delay_unit_5.forward.t0 variable_delay_unit_5.in.t3 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X26 VSS.t89 variable_delay_unit_4.tristate_inverter_1.en.t2 a_14288_352# VSS.t88 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X27 VSS.t30 en_1.t2 a_4562_352# VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X28 variable_delay_unit_0.tristate_inverter_1.en.t0 en_0.t2 VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X29 VSS.t40 variable_delay_unit_3.tristate_inverter_1.en.t2 a_11340_352# VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X30 variable_delay_unit_5.in.t1 variable_delay_unit_4.in.t2 VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X31 VDD.t18 variable_delay_unit_4.tristate_inverter_1.en.t3 a_13406_772# VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X32 variable_delay_unit_3.out variable_delay_unit_4.in.t3 a_10458_772# VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X33 out.t3 variable_delay_unit_1.in.t3 a_1614_352# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X34 VDD.t20 en_2.t1 a_8392_772# VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X35 variable_delay_unit_5.in.t0 variable_delay_unit_4.in.t4 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X36 VSS.t53 en_4.t1 a_13406_352# VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X37 variable_delay_unit_3.out variable_delay_unit_4.in.t5 a_10458_352# VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X38 a_2496_772# variable_delay_unit_1.out out.t1 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X39 VDD.t77 VDD.t75 a_17236_772# VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X40 VDD.t66 variable_delay_unit_3.tristate_inverter_1.en.t3 a_10458_772# VDD.t65 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X41 VSS.t69 variable_delay_unit_2.tristate_inverter_1.en.t4 a_8392_352# VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X42 VSS.t83 variable_delay_unit_5.tristate_inverter_1.en.t4 a_17236_352# VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X43 variable_delay_unit_2.out variable_delay_unit_3.in.t4 a_7510_772# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X44 a_2496_352# variable_delay_unit_1.out out.t0 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X45 VSS.t55 en_3.t1 a_10458_352# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X46 VDD.t30 en_4.t2 a_14288_772# VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X47 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t3 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X48 variable_delay_unit_2.out variable_delay_unit_3.in.t5 a_7510_352# VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X49 VSS.t99 variable_delay_unit_4.tristate_inverter_1.en.t4 a_14288_352# VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X50 a_1614_352# en_0.t3 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X51 variable_delay_unit_5.out variable_delay_unit_5.forward.t2 a_16354_772# VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X52 a_5444_772# en_1.t3 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X53 a_8392_772# variable_delay_unit_3.out variable_delay_unit_2.out VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X54 VDD.t84 variable_delay_unit_5.tristate_inverter_1.en.t5 a_16354_772# VDD.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X55 variable_delay_unit_4.out variable_delay_unit_5.in.t4 a_13406_772# VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X56 variable_delay_unit_1.tristate_inverter_1.en.t1 en_1.t4 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X57 variable_delay_unit_5.out variable_delay_unit_5.forward.t3 a_16354_352# VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X58 a_8392_352# variable_delay_unit_3.out variable_delay_unit_2.out VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X59 VSS.t77 VDD.t113 a_16354_352# VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X60 a_5444_352# variable_delay_unit_1.tristate_inverter_1.en.t5 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X61 variable_delay_unit_4.out variable_delay_unit_5.in.t5 a_13406_352# VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X62 a_5444_772# variable_delay_unit_2.out variable_delay_unit_1.out VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X63 variable_delay_unit_1.tristate_inverter_1.en.t0 en_1.t5 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X64 a_2496_772# en_0.t4 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X65 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en.t5 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X66 a_5444_352# variable_delay_unit_2.out variable_delay_unit_1.out VSS.t101 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X67 a_2496_352# variable_delay_unit_0.tristate_inverter_1.en.t4 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X68 a_7510_352# en_2.t2 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X69 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t6 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X70 a_14288_772# variable_delay_unit_5.out variable_delay_unit_4.out VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X71 a_11340_772# en_3.t2 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X72 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en.t5 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X73 variable_delay_unit_3.tristate_inverter_1.en.t1 en_3.t3 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X74 a_11340_772# variable_delay_unit_4.out variable_delay_unit_3.out VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X75 a_14288_352# variable_delay_unit_5.out variable_delay_unit_4.out VSS.t92 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X76 a_4562_352# en_1.t6 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X77 a_11340_352# variable_delay_unit_3.tristate_inverter_1.en.t4 VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X78 variable_delay_unit_3.tristate_inverter_1.en.t0 en_3.t4 VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X79 a_1614_352# en_0.t5 VSS.t108 VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X80 variable_delay_unit_1.in.t0 in.t0 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X81 a_11340_352# variable_delay_unit_4.out variable_delay_unit_3.out VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X82 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en.t5 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X83 variable_delay_unit_2.tristate_inverter_1.en.t0 en_2.t3 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X84 a_8392_772# en_2.t4 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X85 variable_delay_unit_1.in.t1 in.t1 VSS.t106 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X86 a_13406_352# en_4.t3 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X87 variable_delay_unit_2.tristate_inverter_1.en.t1 en_2.t5 VSS.t87 VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X88 a_17236_772# VDD.t72 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X89 a_8392_352# variable_delay_unit_2.tristate_inverter_1.en.t6 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X90 a_10458_772# variable_delay_unit_3.tristate_inverter_1.en.t5 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X91 variable_delay_unit_5.tristate_inverter_1.en.t1 VDD.t69 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X92 a_17236_352# variable_delay_unit_5.tristate_inverter_1.en.t6 VSS.t81 VSS.t80 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X93 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en.t7 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X94 a_10458_352# en_3.t5 VSS.t42 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X95 variable_delay_unit_5.tristate_inverter_1.en.t0 VDD.t114 VSS.t75 VSS.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X96 a_17236_772# VSS.t109 variable_delay_unit_5.out VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X97 a_14288_772# en_4.t4 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X98 a_7510_352# en_2.t6 VSS.t22 VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X99 variable_delay_unit_4.tristate_inverter_1.en.t1 en_4.t5 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X100 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en.t7 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X101 a_17236_352# VSS.t15 variable_delay_unit_5.out VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X102 a_14288_352# variable_delay_unit_4.tristate_inverter_1.en.t6 VSS.t57 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X103 variable_delay_unit_4.tristate_inverter_1.en.t0 en_4.t6 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X104 a_16354_772# variable_delay_unit_5.tristate_inverter_1.en.t7 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X105 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en.t7 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X106 a_4562_352# en_1.t7 VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X107 a_16354_352# VDD.t115 VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X108 a_13406_352# en_4.t7 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X109 VDD.t35 en_0.t6 a_2496_772# VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X110 variable_delay_unit_2.in.t0 variable_delay_unit_1.in.t4 VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X111 a_10458_772# variable_delay_unit_3.tristate_inverter_1.en.t6 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X112 variable_delay_unit_2.in.t1 variable_delay_unit_1.in.t5 VSS.t94 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X113 VSS.t97 variable_delay_unit_0.tristate_inverter_1.en.t6 a_2496_352# VSS.t96 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X114 a_10458_352# en_3.t6 VSS.t38 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X115 VDD.t48 variable_delay_unit_0.tristate_inverter_1.en.t7 a_1614_772# VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X116 VDD.t16 en_3.t7 a_11340_772# VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X117 VSS.t34 en_0.t7 a_1614_352# VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X118 VSS.t91 variable_delay_unit_3.tristate_inverter_1.en.t7 a_11340_352# VSS.t90 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X119 VDD.t88 en_2.t7 a_8392_772# VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
R0 variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_unit_5.tristate_inverter_1.en.t7 628.097
R1 variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_unit_5.tristate_inverter_1.en.t2 622.766
R2 variable_delay_unit_5.tristate_inverter_1.en.n3 variable_delay_unit_5.tristate_inverter_1.en.t5 523.774
R3 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t3 304.647
R4 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t4 304.647
R5 variable_delay_unit_5.tristate_inverter_1.en.n0 variable_delay_unit_5.tristate_inverter_1.en.t6 202.44
R6 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n0 168.969
R7 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n4 166.147
R8 variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_unit_5.tristate_inverter_1.en.t1 84.7557
R9 variable_delay_unit_5.tristate_inverter_1.en.n1 variable_delay_unit_5.tristate_inverter_1.en.t0 84.1197
R10 variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_unit_5.tristate_inverter_1.en.n1 12.6535
R11 variable_delay_unit_5.tristate_inverter_1.en.n2 variable_delay_unit_5.tristate_inverter_1.en 5.58443
R12 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en.n2 4.59003
R13 variable_delay_unit_5.tristate_inverter_1.en.n4 variable_delay_unit_5.tristate_inverter_1.en.n3 1.09595
R14 VDD.n298 VDD.n264 1689.71
R15 VDD.n269 VDD.n264 1689.71
R16 VDD.n262 VDD.n261 1689.71
R17 VDD.n301 VDD.n261 1689.71
R18 VDD.n238 VDD.n13 1689.71
R19 VDD.n238 VDD.n14 1689.71
R20 VDD.n20 VDD.n15 1689.71
R21 VDD.n234 VDD.n15 1689.71
R22 VDD.n210 VDD.n35 1689.71
R23 VDD.n210 VDD.n36 1689.71
R24 VDD.n42 VDD.n37 1689.71
R25 VDD.n206 VDD.n37 1689.71
R26 VDD.n182 VDD.n57 1689.71
R27 VDD.n182 VDD.n58 1689.71
R28 VDD.n64 VDD.n59 1689.71
R29 VDD.n178 VDD.n59 1689.71
R30 VDD.n154 VDD.n79 1689.71
R31 VDD.n154 VDD.n80 1689.71
R32 VDD.n86 VDD.n81 1689.71
R33 VDD.n150 VDD.n81 1689.71
R34 VDD.n118 VDD.n101 1689.71
R35 VDD.n118 VDD.n102 1689.71
R36 VDD.n108 VDD.n103 1689.71
R37 VDD.n114 VDD.n103 1689.71
R38 VDD.n132 VDD.n91 1307.92
R39 VDD.n128 VDD.n92 1307.92
R40 VDD.n168 VDD.n69 1307.92
R41 VDD.n164 VDD.n70 1307.92
R42 VDD.n196 VDD.n47 1307.92
R43 VDD.n192 VDD.n48 1307.92
R44 VDD.n224 VDD.n25 1307.92
R45 VDD.n220 VDD.n26 1307.92
R46 VDD.n252 VDD.n3 1307.92
R47 VDD.n248 VDD.n4 1307.92
R48 VDD.n281 VDD.n277 1307.92
R49 VDD.n274 VDD.n273 1307.92
R50 VDD.n138 VDD.t75 628.097
R51 VDD.n139 VDD.t78 622.766
R52 VDD.n142 VDD.t69 543.053
R53 VDD.n138 VDD.t72 523.774
R54 VDD.n300 VDD.n299 332.803
R55 VDD.n236 VDD.n235 332.803
R56 VDD.n208 VDD.n207 332.803
R57 VDD.n180 VDD.n179 332.803
R58 VDD.n152 VDD.n151 332.803
R59 VDD.n116 VDD.n115 332.803
R60 VDD.n137 VDD.t115 304.647
R61 VDD.n137 VDD.t112 304.647
R62 VDD.n142 VDD.t114 221.72
R63 VDD.n143 VDD.n142 219.526
R64 VDD.n137 VDD.t113 202.44
R65 VDD.n297 VDD.n265 180.236
R66 VDD.n270 VDD.n265 180.236
R67 VDD.n303 VDD.n302 180.236
R68 VDD.n303 VDD.n257 180.236
R69 VDD.n239 VDD.n12 180.236
R70 VDD.n239 VDD.n8 180.236
R71 VDD.n233 VDD.n16 180.236
R72 VDD.n21 VDD.n16 180.236
R73 VDD.n211 VDD.n34 180.236
R74 VDD.n211 VDD.n30 180.236
R75 VDD.n205 VDD.n38 180.236
R76 VDD.n43 VDD.n38 180.236
R77 VDD.n183 VDD.n56 180.236
R78 VDD.n183 VDD.n52 180.236
R79 VDD.n177 VDD.n60 180.236
R80 VDD.n65 VDD.n60 180.236
R81 VDD.n155 VDD.n78 180.236
R82 VDD.n155 VDD.n74 180.236
R83 VDD.n149 VDD.n82 180.236
R84 VDD.n87 VDD.n82 180.236
R85 VDD.n119 VDD.n100 180.236
R86 VDD.n119 VDD.n96 180.236
R87 VDD.n113 VDD.n104 180.236
R88 VDD.n109 VDD.n104 180.236
R89 VDD.n131 VDD.n88 175.123
R90 VDD.n95 VDD.n94 175.123
R91 VDD.n167 VDD.n66 175.123
R92 VDD.n73 VDD.n72 175.123
R93 VDD.n195 VDD.n44 175.123
R94 VDD.n51 VDD.n50 175.123
R95 VDD.n223 VDD.n22 175.123
R96 VDD.n29 VDD.n28 175.123
R97 VDD.n251 VDD.n0 175.123
R98 VDD.n7 VDD.n6 175.123
R99 VDD.n284 VDD.n283 175.123
R100 VDD.n279 VDD.n271 175.123
R101 VDD VDD.n137 168.969
R102 VDD VDD.n139 166.147
R103 VDD.t49 VDD.n262 163.724
R104 VDD.n269 VDD.t5 163.724
R105 VDD.n20 VDD.t53 163.724
R106 VDD.t45 VDD.n14 163.724
R107 VDD.n42 VDD.t19 163.724
R108 VDD.t91 VDD.n36 163.724
R109 VDD.n64 VDD.t51 163.724
R110 VDD.t97 VDD.n58 163.724
R111 VDD.n86 VDD.t29 163.724
R112 VDD.t7 VDD.n80 163.724
R113 VDD.n108 VDD.t76 163.724
R114 VDD.t81 VDD.n102 163.724
R115 VDD.n129 VDD.t95 160.923
R116 VDD.t70 VDD.n130 160.923
R117 VDD.n165 VDD.t109 160.923
R118 VDD.t1 VDD.n166 160.923
R119 VDD.n193 VDD.t3 160.923
R120 VDD.t58 VDD.n194 160.923
R121 VDD.n221 VDD.t39 160.923
R122 VDD.t32 VDD.n222 160.923
R123 VDD.n249 VDD.t101 160.923
R124 VDD.t11 VDD.n250 160.923
R125 VDD.n280 VDD.t89 160.923
R126 VDD.t25 VDD.n282 160.923
R127 VDD.n300 VDD.t67 145.224
R128 VDD.n299 VDD.t60 145.224
R129 VDD.n235 VDD.t106 145.224
R130 VDD.t68 VDD.n236 145.224
R131 VDD.n207 VDD.t104 145.224
R132 VDD.t0 VDD.n208 145.224
R133 VDD.n179 VDD.t105 145.224
R134 VDD.t111 VDD.n180 145.224
R135 VDD.n151 VDD.t103 145.224
R136 VDD.t55 VDD.n152 145.224
R137 VDD.n115 VDD.t36 145.224
R138 VDD.t31 VDD.n116 145.224
R139 VDD.n133 VDD.n90 139.512
R140 VDD.n133 VDD.n88 139.512
R141 VDD.n127 VDD.n93 139.512
R142 VDD.n95 VDD.n93 139.512
R143 VDD.n169 VDD.n68 139.512
R144 VDD.n169 VDD.n66 139.512
R145 VDD.n163 VDD.n71 139.512
R146 VDD.n73 VDD.n71 139.512
R147 VDD.n197 VDD.n46 139.512
R148 VDD.n197 VDD.n44 139.512
R149 VDD.n191 VDD.n49 139.512
R150 VDD.n51 VDD.n49 139.512
R151 VDD.n225 VDD.n24 139.512
R152 VDD.n225 VDD.n22 139.512
R153 VDD.n219 VDD.n27 139.512
R154 VDD.n29 VDD.n27 139.512
R155 VDD.n253 VDD.n2 139.512
R156 VDD.n253 VDD.n0 139.512
R157 VDD.n247 VDD.n5 139.512
R158 VDD.n7 VDD.n5 139.512
R159 VDD.n285 VDD.n275 139.512
R160 VDD.n285 VDD.n284 139.512
R161 VDD.n290 VDD.n289 139.512
R162 VDD.n290 VDD.n271 139.512
R163 VDD.n130 VDD.n129 119.861
R164 VDD.n166 VDD.n165 119.861
R165 VDD.n194 VDD.n193 119.861
R166 VDD.n222 VDD.n221 119.861
R167 VDD.n250 VDD.n249 119.861
R168 VDD.n282 VDD.n280 119.861
R169 VDD.t27 VDD.t49 88.7478
R170 VDD.t67 VDD.t34 88.7478
R171 VDD.t99 VDD.t60 88.7478
R172 VDD.t5 VDD.t47 88.7478
R173 VDD.t53 VDD.t13 88.7478
R174 VDD.t23 VDD.t106 88.7478
R175 VDD.t21 VDD.t68 88.7478
R176 VDD.t107 VDD.t45 88.7478
R177 VDD.t19 VDD.t41 88.7478
R178 VDD.t87 VDD.t104 88.7478
R179 VDD.t37 VDD.t0 88.7478
R180 VDD.t93 VDD.t91 88.7478
R181 VDD.t51 VDD.t9 88.7478
R182 VDD.t15 VDD.t105 88.7478
R183 VDD.t63 VDD.t111 88.7478
R184 VDD.t65 VDD.t97 88.7478
R185 VDD.t29 VDD.t43 88.7478
R186 VDD.t56 VDD.t103 88.7478
R187 VDD.t61 VDD.t55 88.7478
R188 VDD.t17 VDD.t7 88.7478
R189 VDD.t76 VDD.t73 88.7478
R190 VDD.t79 VDD.t36 88.7478
R191 VDD.t85 VDD.t31 88.7478
R192 VDD.t83 VDD.t81 88.7478
R193 VDD.n135 VDD.t71 84.7934
R194 VDD.n125 VDD.t96 84.7934
R195 VDD.n171 VDD.t2 84.7934
R196 VDD.n161 VDD.t110 84.7934
R197 VDD.n199 VDD.t59 84.7934
R198 VDD.n189 VDD.t4 84.7934
R199 VDD.n227 VDD.t33 84.7934
R200 VDD.n217 VDD.t40 84.7934
R201 VDD.n255 VDD.t12 84.7934
R202 VDD.n245 VDD.t102 84.7934
R203 VDD.n276 VDD.t26 84.7934
R204 VDD.n272 VDD.t90 84.7934
R205 VDD.n267 VDD.n266 84.7744
R206 VDD.n259 VDD.n258 84.7744
R207 VDD.n10 VDD.n9 84.7744
R208 VDD.n18 VDD.n17 84.7744
R209 VDD.n32 VDD.n31 84.7744
R210 VDD.n40 VDD.n39 84.7744
R211 VDD.n54 VDD.n53 84.7744
R212 VDD.n62 VDD.n61 84.7744
R213 VDD.n76 VDD.n75 84.7744
R214 VDD.n84 VDD.n83 84.7744
R215 VDD.n98 VDD.n97 84.7744
R216 VDD.n106 VDD.n105 84.7744
R217 VDD.n267 VDD.t6 83.8097
R218 VDD.n259 VDD.t50 83.8097
R219 VDD.n10 VDD.t46 83.8097
R220 VDD.n18 VDD.t54 83.8097
R221 VDD.n32 VDD.t92 83.8097
R222 VDD.n40 VDD.t20 83.8097
R223 VDD.n54 VDD.t98 83.8097
R224 VDD.n62 VDD.t52 83.8097
R225 VDD.n76 VDD.t8 83.8097
R226 VDD.n84 VDD.t30 83.8097
R227 VDD.n98 VDD.t82 83.8097
R228 VDD.n106 VDD.t77 83.8097
R229 VDD.n133 VDD.n132 46.2505
R230 VDD.n93 VDD.n92 46.2505
R231 VDD.n169 VDD.n168 46.2505
R232 VDD.n71 VDD.n70 46.2505
R233 VDD.n197 VDD.n196 46.2505
R234 VDD.n49 VDD.n48 46.2505
R235 VDD.n225 VDD.n224 46.2505
R236 VDD.n27 VDD.n26 46.2505
R237 VDD.n253 VDD.n252 46.2505
R238 VDD.n5 VDD.n4 46.2505
R239 VDD.n285 VDD.n277 46.2505
R240 VDD.n290 VDD.n273 46.2505
R241 VDD.n263 VDD.t27 44.3742
R242 VDD.t34 VDD.n263 44.3742
R243 VDD.n268 VDD.t99 44.3742
R244 VDD.t47 VDD.n268 44.3742
R245 VDD.t13 VDD.n19 44.3742
R246 VDD.n19 VDD.t23 44.3742
R247 VDD.n237 VDD.t21 44.3742
R248 VDD.n237 VDD.t107 44.3742
R249 VDD.t41 VDD.n41 44.3742
R250 VDD.n41 VDD.t87 44.3742
R251 VDD.n209 VDD.t37 44.3742
R252 VDD.n209 VDD.t93 44.3742
R253 VDD.t9 VDD.n63 44.3742
R254 VDD.n63 VDD.t15 44.3742
R255 VDD.n181 VDD.t63 44.3742
R256 VDD.n181 VDD.t65 44.3742
R257 VDD.t43 VDD.n85 44.3742
R258 VDD.n85 VDD.t56 44.3742
R259 VDD.n153 VDD.t61 44.3742
R260 VDD.n153 VDD.t17 44.3742
R261 VDD.t73 VDD.n107 44.3742
R262 VDD.n107 VDD.t79 44.3742
R263 VDD.n117 VDD.t85 44.3742
R264 VDD.n117 VDD.t83 44.3742
R265 VDD.n132 VDD.n131 39.3924
R266 VDD.n94 VDD.n92 39.3924
R267 VDD.n168 VDD.n167 39.3924
R268 VDD.n72 VDD.n70 39.3924
R269 VDD.n196 VDD.n195 39.3924
R270 VDD.n50 VDD.n48 39.3924
R271 VDD.n224 VDD.n223 39.3924
R272 VDD.n28 VDD.n26 39.3924
R273 VDD.n252 VDD.n251 39.3924
R274 VDD.n6 VDD.n4 39.3924
R275 VDD.n283 VDD.n277 39.3924
R276 VDD.n279 VDD.n273 39.3924
R277 VDD.n265 VDD.n264 23.1255
R278 VDD.n268 VDD.n264 23.1255
R279 VDD.n303 VDD.n261 23.1255
R280 VDD.n263 VDD.n261 23.1255
R281 VDD.n239 VDD.n238 23.1255
R282 VDD.n238 VDD.n237 23.1255
R283 VDD.n16 VDD.n15 23.1255
R284 VDD.n19 VDD.n15 23.1255
R285 VDD.n211 VDD.n210 23.1255
R286 VDD.n210 VDD.n209 23.1255
R287 VDD.n38 VDD.n37 23.1255
R288 VDD.n41 VDD.n37 23.1255
R289 VDD.n183 VDD.n182 23.1255
R290 VDD.n182 VDD.n181 23.1255
R291 VDD.n60 VDD.n59 23.1255
R292 VDD.n63 VDD.n59 23.1255
R293 VDD.n155 VDD.n154 23.1255
R294 VDD.n154 VDD.n153 23.1255
R295 VDD.n82 VDD.n81 23.1255
R296 VDD.n85 VDD.n81 23.1255
R297 VDD.n119 VDD.n118 23.1255
R298 VDD.n118 VDD.n117 23.1255
R299 VDD.n104 VDD.n103 23.1255
R300 VDD.n107 VDD.n103 23.1255
R301 VDD.n91 VDD.n90 20.5561
R302 VDD.n130 VDD.n91 20.5561
R303 VDD.n128 VDD.n127 20.5561
R304 VDD.n129 VDD.n128 20.5561
R305 VDD.n69 VDD.n68 20.5561
R306 VDD.n166 VDD.n69 20.5561
R307 VDD.n164 VDD.n163 20.5561
R308 VDD.n165 VDD.n164 20.5561
R309 VDD.n47 VDD.n46 20.5561
R310 VDD.n194 VDD.n47 20.5561
R311 VDD.n192 VDD.n191 20.5561
R312 VDD.n193 VDD.n192 20.5561
R313 VDD.n25 VDD.n24 20.5561
R314 VDD.n222 VDD.n25 20.5561
R315 VDD.n220 VDD.n219 20.5561
R316 VDD.n221 VDD.n220 20.5561
R317 VDD.n3 VDD.n2 20.5561
R318 VDD.n250 VDD.n3 20.5561
R319 VDD.n248 VDD.n247 20.5561
R320 VDD.n249 VDD.n248 20.5561
R321 VDD.n281 VDD.n275 20.5561
R322 VDD.n282 VDD.n281 20.5561
R323 VDD.n289 VDD.n274 20.5561
R324 VDD.n280 VDD.n274 20.5561
R325 VDD.n270 VDD.n269 18.5005
R326 VDD.n298 VDD.n297 18.5005
R327 VDD.n299 VDD.n298 18.5005
R328 VDD.n302 VDD.n301 18.5005
R329 VDD.n301 VDD.n300 18.5005
R330 VDD.n262 VDD.n257 18.5005
R331 VDD.n14 VDD.n8 18.5005
R332 VDD.n13 VDD.n12 18.5005
R333 VDD.n236 VDD.n13 18.5005
R334 VDD.n234 VDD.n233 18.5005
R335 VDD.n235 VDD.n234 18.5005
R336 VDD.n21 VDD.n20 18.5005
R337 VDD.n36 VDD.n30 18.5005
R338 VDD.n35 VDD.n34 18.5005
R339 VDD.n208 VDD.n35 18.5005
R340 VDD.n206 VDD.n205 18.5005
R341 VDD.n207 VDD.n206 18.5005
R342 VDD.n43 VDD.n42 18.5005
R343 VDD.n58 VDD.n52 18.5005
R344 VDD.n57 VDD.n56 18.5005
R345 VDD.n180 VDD.n57 18.5005
R346 VDD.n178 VDD.n177 18.5005
R347 VDD.n179 VDD.n178 18.5005
R348 VDD.n65 VDD.n64 18.5005
R349 VDD.n80 VDD.n74 18.5005
R350 VDD.n79 VDD.n78 18.5005
R351 VDD.n152 VDD.n79 18.5005
R352 VDD.n150 VDD.n149 18.5005
R353 VDD.n151 VDD.n150 18.5005
R354 VDD.n87 VDD.n86 18.5005
R355 VDD.n102 VDD.n96 18.5005
R356 VDD.n101 VDD.n100 18.5005
R357 VDD.n116 VDD.n101 18.5005
R358 VDD.n114 VDD.n113 18.5005
R359 VDD.n115 VDD.n114 18.5005
R360 VDD.n109 VDD.n108 18.5005
R361 VDD.n266 VDD.t100 9.52217
R362 VDD.n266 VDD.t48 9.52217
R363 VDD.n258 VDD.t28 9.52217
R364 VDD.n258 VDD.t35 9.52217
R365 VDD.n9 VDD.t22 9.52217
R366 VDD.n9 VDD.t108 9.52217
R367 VDD.n17 VDD.t14 9.52217
R368 VDD.n17 VDD.t24 9.52217
R369 VDD.n31 VDD.t38 9.52217
R370 VDD.n31 VDD.t94 9.52217
R371 VDD.n39 VDD.t42 9.52217
R372 VDD.n39 VDD.t88 9.52217
R373 VDD.n53 VDD.t64 9.52217
R374 VDD.n53 VDD.t66 9.52217
R375 VDD.n61 VDD.t10 9.52217
R376 VDD.n61 VDD.t16 9.52217
R377 VDD.n75 VDD.t62 9.52217
R378 VDD.n75 VDD.t18 9.52217
R379 VDD.n83 VDD.t44 9.52217
R380 VDD.n83 VDD.t57 9.52217
R381 VDD.n97 VDD.t86 9.52217
R382 VDD.n97 VDD.t84 9.52217
R383 VDD.n105 VDD.t74 9.52217
R384 VDD.n105 VDD.t80 9.52217
R385 VDD.n94 VDD.t95 5.4667
R386 VDD.n131 VDD.t70 5.4667
R387 VDD.n72 VDD.t109 5.4667
R388 VDD.n167 VDD.t1 5.4667
R389 VDD.n50 VDD.t3 5.4667
R390 VDD.n195 VDD.t58 5.4667
R391 VDD.n28 VDD.t39 5.4667
R392 VDD.n223 VDD.t32 5.4667
R393 VDD.n6 VDD.t101 5.4667
R394 VDD.n251 VDD.t11 5.4667
R395 VDD.t89 VDD.n279 5.4667
R396 VDD.n283 VDD.t25 5.4667
R397 VDD.n141 VDD.n140 3.26479
R398 VDD.n124 VDD.n93 2.3255
R399 VDD.n134 VDD.n133 2.3255
R400 VDD.n160 VDD.n71 2.3255
R401 VDD.n170 VDD.n169 2.3255
R402 VDD.n188 VDD.n49 2.3255
R403 VDD.n198 VDD.n197 2.3255
R404 VDD.n216 VDD.n27 2.3255
R405 VDD.n226 VDD.n225 2.3255
R406 VDD.n244 VDD.n5 2.3255
R407 VDD.n254 VDD.n253 2.3255
R408 VDD.n291 VDD.n290 2.3255
R409 VDD.n286 VDD.n285 2.3255
R410 VDD.n144 VDD.n143 2.2505
R411 VDD.n127 VDD.n126 2.04321
R412 VDD.n136 VDD.n88 2.04321
R413 VDD.n90 VDD.n89 2.04321
R414 VDD.n123 VDD.n95 2.04321
R415 VDD.n163 VDD.n162 2.04321
R416 VDD.n172 VDD.n66 2.04321
R417 VDD.n68 VDD.n67 2.04321
R418 VDD.n159 VDD.n73 2.04321
R419 VDD.n191 VDD.n190 2.04321
R420 VDD.n200 VDD.n44 2.04321
R421 VDD.n46 VDD.n45 2.04321
R422 VDD.n187 VDD.n51 2.04321
R423 VDD.n219 VDD.n218 2.04321
R424 VDD.n228 VDD.n22 2.04321
R425 VDD.n24 VDD.n23 2.04321
R426 VDD.n215 VDD.n29 2.04321
R427 VDD.n247 VDD.n246 2.04321
R428 VDD.n256 VDD.n0 2.04321
R429 VDD.n2 VDD.n1 2.04321
R430 VDD.n243 VDD.n7 2.04321
R431 VDD.n289 VDD.n288 2.04321
R432 VDD.n284 VDD.n278 2.04321
R433 VDD.n287 VDD.n275 2.04321
R434 VDD.n292 VDD.n271 2.04321
R435 VDD VDD.n109 1.97234
R436 VDD.n302 VDD.n260 1.96583
R437 VDD.n293 VDD.n270 1.96583
R438 VDD.n297 VDD.n296 1.96583
R439 VDD.n306 VDD.n257 1.96583
R440 VDD.n233 VDD.n232 1.96583
R441 VDD.n242 VDD.n8 1.96583
R442 VDD.n12 VDD.n11 1.96583
R443 VDD.n229 VDD.n21 1.96583
R444 VDD.n205 VDD.n204 1.96583
R445 VDD.n214 VDD.n30 1.96583
R446 VDD.n34 VDD.n33 1.96583
R447 VDD.n201 VDD.n43 1.96583
R448 VDD.n177 VDD.n176 1.96583
R449 VDD.n186 VDD.n52 1.96583
R450 VDD.n56 VDD.n55 1.96583
R451 VDD.n173 VDD.n65 1.96583
R452 VDD.n149 VDD.n148 1.96583
R453 VDD.n158 VDD.n74 1.96583
R454 VDD.n78 VDD.n77 1.96583
R455 VDD.n145 VDD.n87 1.96583
R456 VDD.n113 VDD.n112 1.96583
R457 VDD.n122 VDD.n96 1.96583
R458 VDD.n100 VDD.n99 1.96583
R459 VDD.n140 VDD 1.40175
R460 VDD.n111 VDD.n104 1.32907
R461 VDD.n120 VDD.n119 1.32907
R462 VDD.n147 VDD.n82 1.32907
R463 VDD.n156 VDD.n155 1.32907
R464 VDD.n175 VDD.n60 1.32907
R465 VDD.n184 VDD.n183 1.32907
R466 VDD.n203 VDD.n38 1.32907
R467 VDD.n212 VDD.n211 1.32907
R468 VDD.n231 VDD.n16 1.32907
R469 VDD.n240 VDD.n239 1.32907
R470 VDD.n304 VDD.n303 1.32907
R471 VDD.n295 VDD.n265 1.32907
R472 VDD.n294 VDD.n267 1.21789
R473 VDD.n305 VDD.n259 1.21789
R474 VDD.n241 VDD.n10 1.21789
R475 VDD.n230 VDD.n18 1.21789
R476 VDD.n213 VDD.n32 1.21789
R477 VDD.n202 VDD.n40 1.21789
R478 VDD.n185 VDD.n54 1.21789
R479 VDD.n174 VDD.n62 1.21789
R480 VDD.n157 VDD.n76 1.21789
R481 VDD.n146 VDD.n84 1.21789
R482 VDD.n121 VDD.n98 1.21789
R483 VDD.n110 VDD.n106 1.21789
R484 VDD.n139 VDD.n138 1.09595
R485 VDD.n143 VDD.n141 0.738
R486 VDD VDD.n172 0.568208
R487 VDD VDD.n200 0.568208
R488 VDD VDD.n228 0.568208
R489 VDD VDD.n256 0.568208
R490 VDD.n278 VDD 0.492688
R491 VDD.n140 VDD 0.443357
R492 VDD.n123 VDD 0.432792
R493 VDD.n159 VDD 0.432792
R494 VDD.n187 VDD 0.432792
R495 VDD.n215 VDD 0.432792
R496 VDD.n243 VDD 0.432792
R497 VDD VDD.n292 0.432792
R498 VDD.n112 VDD.n99 0.430188
R499 VDD.n148 VDD.n77 0.430188
R500 VDD.n176 VDD.n55 0.430188
R501 VDD.n204 VDD.n33 0.430188
R502 VDD.n232 VDD.n11 0.430188
R503 VDD.n296 VDD.n260 0.430188
R504 VDD VDD.n144 0.389823
R505 VDD.n112 VDD.n111 0.359875
R506 VDD.n120 VDD.n99 0.359875
R507 VDD.n148 VDD.n147 0.359875
R508 VDD.n156 VDD.n77 0.359875
R509 VDD.n176 VDD.n175 0.359875
R510 VDD.n184 VDD.n55 0.359875
R511 VDD.n204 VDD.n203 0.359875
R512 VDD.n212 VDD.n33 0.359875
R513 VDD.n232 VDD.n231 0.359875
R514 VDD.n240 VDD.n11 0.359875
R515 VDD.n304 VDD.n260 0.359875
R516 VDD.n296 VDD.n295 0.359875
R517 VDD.n111 VDD.n110 0.229667
R518 VDD.n121 VDD.n120 0.229667
R519 VDD.n147 VDD.n146 0.229667
R520 VDD.n157 VDD.n156 0.229667
R521 VDD.n175 VDD.n174 0.229667
R522 VDD.n185 VDD.n184 0.229667
R523 VDD.n203 VDD.n202 0.229667
R524 VDD.n213 VDD.n212 0.229667
R525 VDD.n231 VDD.n230 0.229667
R526 VDD.n241 VDD.n240 0.229667
R527 VDD.n305 VDD.n304 0.229667
R528 VDD.n295 VDD.n294 0.229667
R529 VDD.n124 VDD.n123 0.189302
R530 VDD.n134 VDD.n89 0.189302
R531 VDD.n160 VDD.n159 0.189302
R532 VDD.n170 VDD.n67 0.189302
R533 VDD.n188 VDD.n187 0.189302
R534 VDD.n198 VDD.n45 0.189302
R535 VDD.n216 VDD.n215 0.189302
R536 VDD.n226 VDD.n23 0.189302
R537 VDD.n244 VDD.n243 0.189302
R538 VDD.n254 VDD.n1 0.189302
R539 VDD.n292 VDD.n291 0.189302
R540 VDD.n287 VDD.n286 0.189302
R541 VDD.n144 VDD.n136 0.178885
R542 VDD.n126 VDD.n89 0.141125
R543 VDD.n162 VDD.n67 0.141125
R544 VDD.n190 VDD.n45 0.141125
R545 VDD.n218 VDD.n23 0.141125
R546 VDD.n246 VDD.n1 0.141125
R547 VDD.n288 VDD.n287 0.141125
R548 VDD.n126 VDD.n125 0.13201
R549 VDD.n136 VDD.n135 0.13201
R550 VDD.n162 VDD.n161 0.13201
R551 VDD.n172 VDD.n171 0.13201
R552 VDD.n190 VDD.n189 0.13201
R553 VDD.n200 VDD.n199 0.13201
R554 VDD.n218 VDD.n217 0.13201
R555 VDD.n228 VDD.n227 0.13201
R556 VDD.n246 VDD.n245 0.13201
R557 VDD.n256 VDD.n255 0.13201
R558 VDD.n288 VDD.n272 0.13201
R559 VDD.n278 VDD.n276 0.13201
R560 VDD.n122 VDD.n121 0.130708
R561 VDD.n158 VDD.n157 0.130708
R562 VDD.n186 VDD.n185 0.130708
R563 VDD.n214 VDD.n213 0.130708
R564 VDD.n242 VDD.n241 0.130708
R565 VDD.n294 VDD.n293 0.130708
R566 VDD.n110 VDD 0.124198
R567 VDD.n146 VDD 0.124198
R568 VDD.n174 VDD 0.124198
R569 VDD.n202 VDD 0.124198
R570 VDD.n230 VDD 0.124198
R571 VDD VDD.n305 0.124198
R572 VDD VDD.n122 0.0695104
R573 VDD.n145 VDD 0.0695104
R574 VDD VDD.n158 0.0695104
R575 VDD.n173 VDD 0.0695104
R576 VDD VDD.n186 0.0695104
R577 VDD.n201 VDD 0.0695104
R578 VDD VDD.n214 0.0695104
R579 VDD.n229 VDD 0.0695104
R580 VDD VDD.n242 0.0695104
R581 VDD VDD.n306 0.0695104
R582 VDD.n293 VDD 0.0695104
R583 VDD.n141 VDD 0.063
R584 VDD.n125 VDD.n124 0.0577917
R585 VDD.n135 VDD.n134 0.0577917
R586 VDD.n161 VDD.n160 0.0577917
R587 VDD.n171 VDD.n170 0.0577917
R588 VDD.n189 VDD.n188 0.0577917
R589 VDD.n199 VDD.n198 0.0577917
R590 VDD.n217 VDD.n216 0.0577917
R591 VDD.n227 VDD.n226 0.0577917
R592 VDD.n245 VDD.n244 0.0577917
R593 VDD.n255 VDD.n254 0.0577917
R594 VDD.n291 VDD.n272 0.0577917
R595 VDD.n286 VDD.n276 0.0577917
R596 VDD VDD.n145 0.00701042
R597 VDD VDD.n173 0.00701042
R598 VDD VDD.n201 0.00701042
R599 VDD VDD.n229 0.00701042
R600 VDD.n306 VDD 0.00701042
R601 en_1.n2 en_1.t0 628.097
R602 en_1.n3 en_1.t1 622.766
R603 en_1.n0 en_1.t4 543.053
R604 en_1.n2 en_1.t3 523.774
R605 en_1.n1 en_1.t6 304.647
R606 en_1.n1 en_1.t7 304.647
R607 en_1.n0 en_1.t5 221.72
R608 en_1.n5 en_1.n0 220.263
R609 en_1.n1 en_1.t2 202.44
R610 en_1 en_1.n1 168.969
R611 en_1 en_1.n3 166.147
R612 en_1 en_1.n4 3.15943
R613 en_1.n4 en_1 1.40175
R614 en_1.n3 en_1.n2 1.09595
R615 en_1.n4 en_1 0.443357
R616 en_1.n5 en_1 0.105857
R617 en_1 en_1.n5 0.063
R618 variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_unit_2.tristate_inverter_1.en.t5 628.097
R619 variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_unit_2.tristate_inverter_1.en.t7 622.766
R620 variable_delay_unit_2.tristate_inverter_1.en.n3 variable_delay_unit_2.tristate_inverter_1.en.t3 523.774
R621 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t2 304.647
R622 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t4 304.647
R623 variable_delay_unit_2.tristate_inverter_1.en.n0 variable_delay_unit_2.tristate_inverter_1.en.t6 202.44
R624 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n0 168.969
R625 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n4 166.147
R626 variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_unit_2.tristate_inverter_1.en.t0 84.7557
R627 variable_delay_unit_2.tristate_inverter_1.en.n1 variable_delay_unit_2.tristate_inverter_1.en.t1 84.1197
R628 variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_unit_2.tristate_inverter_1.en.n1 12.6535
R629 variable_delay_unit_2.tristate_inverter_1.en.n2 variable_delay_unit_2.tristate_inverter_1.en 5.58443
R630 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en.n2 4.59003
R631 variable_delay_unit_2.tristate_inverter_1.en.n4 variable_delay_unit_2.tristate_inverter_1.en.n3 1.09595
R632 VSS.n125 VSS.n124 50016.6
R633 VSS.n309 VSS.n308 23663.9
R634 VSS.n212 VSS.n22 23663.9
R635 VSS.n211 VSS.n210 23663.9
R636 VSS.n126 VSS.n52 23663.9
R637 VSS.n317 VSS.n310 23663.9
R638 VSS.n318 VSS.n317 22860.5
R639 VSS.n125 VSS.n81 14239.4
R640 VSS.n147 VSS.n52 14239.4
R641 VSS.n211 VSS.n51 14239.4
R642 VSS.n233 VSS.n22 14239.4
R643 VSS.n309 VSS.n21 14239.4
R644 VSS.n317 VSS.n316 14239.4
R645 VSS.n126 VSS.n125 10823.2
R646 VSS.n210 VSS.n52 10823.2
R647 VSS.n212 VSS.n211 10823.2
R648 VSS.n308 VSS.n22 10823.2
R649 VSS.n310 VSS.n309 10823.2
R650 VSS.n310 VSS.n20 10102.8
R651 VSS.n130 VSS.n126 10102.8
R652 VSS.n210 VSS.n209 10102.8
R653 VSS.n216 VSS.n212 10102.8
R654 VSS.n308 VSS.n307 10102.8
R655 VSS.n112 VSS.n111 2045.07
R656 VSS.n144 VSS.n143 2045.07
R657 VSS.n196 VSS.n195 2045.07
R658 VSS.n230 VSS.n229 2045.07
R659 VSS.n294 VSS.n293 2045.07
R660 VSS.n341 VSS.n340 2045.07
R661 VSS.n342 VSS.n5 1626.7
R662 VSS.n18 VSS.n5 1626.7
R663 VSS.n297 VSS.n291 1626.7
R664 VSS.n297 VSS.n290 1626.7
R665 VSS.n259 VSS.n24 1626.7
R666 VSS.n305 VSS.n24 1626.7
R667 VSS.n236 VSS.n39 1626.7
R668 VSS.n236 VSS.n38 1626.7
R669 VSS.n228 VSS.n40 1626.7
R670 VSS.n214 VSS.n40 1626.7
R671 VSS.n199 VSS.n193 1626.7
R672 VSS.n199 VSS.n192 1626.7
R673 VSS.n173 VSS.n54 1626.7
R674 VSS.n207 VSS.n54 1626.7
R675 VSS.n150 VSS.n69 1626.7
R676 VSS.n150 VSS.n68 1626.7
R677 VSS.n142 VSS.n70 1626.7
R678 VSS.n128 VSS.n70 1626.7
R679 VSS.n115 VSS.n109 1626.7
R680 VSS.n115 VSS.n108 1626.7
R681 VSS.n89 VSS.n82 1626.7
R682 VSS.n123 VSS.n82 1626.7
R683 VSS.n312 VSS.n6 1626.7
R684 VSS.n339 VSS.n6 1626.7
R685 VSS.n209 VSS.n53 1460.78
R686 VSS.n217 VSS.n216 1460.78
R687 VSS.n307 VSS.n23 1460.78
R688 VSS.n272 VSS.n20 1460.78
R689 VSS.n131 VSS.n130 1460.78
R690 VSS.n130 VSS.n129 1437.75
R691 VSS.n209 VSS.n208 1437.75
R692 VSS.n216 VSS.n215 1437.75
R693 VSS.n307 VSS.n306 1437.75
R694 VSS.n20 VSS.n19 1437.75
R695 VSS.n147 VSS.n146 1138.52
R696 VSS.n183 VSS.n51 1138.52
R697 VSS.n233 VSS.n232 1138.52
R698 VSS.n269 VSS.n21 1138.52
R699 VSS.n100 VSS.n81 1138.52
R700 VSS.n316 VSS.n315 1138.52
R701 VSS.n113 VSS.n81 1115.49
R702 VSS.n148 VSS.n147 1115.49
R703 VSS.n197 VSS.n51 1115.49
R704 VSS.n234 VSS.n233 1115.49
R705 VSS.n295 VSS.n21 1115.49
R706 VSS.n316 VSS.n313 1115.49
R707 VSS.n132 VSS.n79 1058.19
R708 VSS.n132 VSS.n78 1058.19
R709 VSS.n102 VSS.n99 1058.19
R710 VSS.n102 VSS.n98 1058.19
R711 VSS.n160 VSS.n60 1058.19
R712 VSS.n145 VSS.n60 1058.19
R713 VSS.n163 VSS.n59 1058.19
R714 VSS.n163 VSS.n58 1058.19
R715 VSS.n185 VSS.n180 1058.19
R716 VSS.n182 VSS.n180 1058.19
R717 VSS.n218 VSS.n49 1058.19
R718 VSS.n218 VSS.n48 1058.19
R719 VSS.n246 VSS.n30 1058.19
R720 VSS.n231 VSS.n30 1058.19
R721 VSS.n249 VSS.n29 1058.19
R722 VSS.n249 VSS.n28 1058.19
R723 VSS.n283 VSS.n266 1058.19
R724 VSS.n268 VSS.n266 1058.19
R725 VSS.n273 VSS.n270 1058.19
R726 VSS.n280 VSS.n270 1058.19
R727 VSS.n319 VSS.n15 1058.19
R728 VSS.n326 VSS.n15 1058.19
R729 VSS.n329 VSS.n13 1058.19
R730 VSS.n314 VSS.n13 1058.19
R731 VSS.n146 VSS.t31 943.788
R732 VSS.n161 VSS.t31 943.788
R733 VSS.t64 VSS.n162 943.788
R734 VSS.t64 VSS.n53 943.788
R735 VSS.t17 VSS.n183 943.788
R736 VSS.n184 VSS.t17 943.788
R737 VSS.t43 VSS.n50 943.788
R738 VSS.t43 VSS.n217 943.788
R739 VSS.n232 VSS.t0 943.788
R740 VSS.n247 VSS.t0 943.788
R741 VSS.t86 VSS.n248 943.788
R742 VSS.t86 VSS.n23 943.788
R743 VSS.t93 VSS.n269 943.788
R744 VSS.n282 VSS.t93 943.788
R745 VSS.n281 VSS.t25 943.788
R746 VSS.n272 VSS.t25 943.788
R747 VSS.t2 VSS.n100 943.788
R748 VSS.t2 VSS.n101 943.788
R749 VSS.t74 VSS.n80 943.788
R750 VSS.t74 VSS.n131 943.788
R751 VSS.n315 VSS.t105 943.788
R752 VSS.n328 VSS.t105 943.788
R753 VSS.n327 VSS.t103 943.788
R754 VSS.n318 VSS.t103 943.788
R755 VSS.n124 VSS.t82 892.394
R756 VSS.n111 VSS.t16 892.394
R757 VSS.t51 VSS.n112 892.394
R758 VSS.t72 VSS.n113 892.394
R759 VSS.n129 VSS.t98 892.394
R760 VSS.n143 VSS.t92 892.394
R761 VSS.t13 VSS.n144 892.394
R762 VSS.t19 VSS.n148 892.394
R763 VSS.n208 VSS.t39 892.394
R764 VSS.n195 VSS.t100 892.394
R765 VSS.t102 VSS.n196 892.394
R766 VSS.t41 VSS.n197 892.394
R767 VSS.n215 VSS.t68 892.394
R768 VSS.n229 VSS.t95 892.394
R769 VSS.t61 VSS.n230 892.394
R770 VSS.t4 VSS.n234 892.394
R771 VSS.n306 VSS.t35 892.394
R772 VSS.n293 VSS.t101 892.394
R773 VSS.t8 VSS.n294 892.394
R774 VSS.t27 VSS.n295 892.394
R775 VSS.n19 VSS.t49 892.394
R776 VSS.n341 VSS.t60 892.394
R777 VSS.n340 VSS.t14 892.394
R778 VSS.n313 VSS.t9 892.394
R779 VSS.n162 VSS.n161 702.96
R780 VSS.n184 VSS.n50 702.96
R781 VSS.n248 VSS.n247 702.96
R782 VSS.n282 VSS.n281 702.96
R783 VSS.n101 VSS.n80 702.96
R784 VSS.n328 VSS.n327 702.96
R785 VSS.n83 VSS.t109 607.409
R786 VSS.t80 VSS.t82 545.352
R787 VSS.t16 VSS.t84 545.352
R788 VSS.t78 VSS.t51 545.352
R789 VSS.t76 VSS.t72 545.352
R790 VSS.t98 VSS.t56 545.352
R791 VSS.t88 VSS.t92 545.352
R792 VSS.t11 VSS.t13 545.352
R793 VSS.t52 VSS.t19 545.352
R794 VSS.t58 VSS.t39 545.352
R795 VSS.t100 VSS.t90 545.352
R796 VSS.t37 VSS.t102 545.352
R797 VSS.t54 VSS.t41 545.352
R798 VSS.t68 VSS.t66 545.352
R799 VSS.t70 VSS.t95 545.352
R800 VSS.t21 VSS.t61 545.352
R801 VSS.t6 VSS.t4 545.352
R802 VSS.t45 VSS.t35 545.352
R803 VSS.t101 VSS.t47 545.352
R804 VSS.t23 VSS.t8 545.352
R805 VSS.t29 VSS.t27 545.352
R806 VSS.t49 VSS.t62 545.352
R807 VSS.t96 VSS.t60 545.352
R808 VSS.t107 VSS.t14 545.352
R809 VSS.t9 VSS.t33 545.352
R810 VSS.n83 VSS.t15 321.423
R811 VSS.n110 VSS.t80 272.676
R812 VSS.t84 VSS.n110 272.676
R813 VSS.n114 VSS.t78 272.676
R814 VSS.n114 VSS.t76 272.676
R815 VSS.t56 VSS.n127 272.676
R816 VSS.n127 VSS.t88 272.676
R817 VSS.n149 VSS.t11 272.676
R818 VSS.n149 VSS.t52 272.676
R819 VSS.n194 VSS.t58 272.676
R820 VSS.t90 VSS.n194 272.676
R821 VSS.n198 VSS.t37 272.676
R822 VSS.n198 VSS.t54 272.676
R823 VSS.t66 VSS.n213 272.676
R824 VSS.n213 VSS.t70 272.676
R825 VSS.n235 VSS.t21 272.676
R826 VSS.n235 VSS.t6 272.676
R827 VSS.n292 VSS.t45 272.676
R828 VSS.t47 VSS.n292 272.676
R829 VSS.n296 VSS.t23 272.676
R830 VSS.n296 VSS.t29 272.676
R831 VSS.t62 VSS.n17 272.676
R832 VSS.n17 VSS.t96 272.676
R833 VSS.n311 VSS.t107 272.676
R834 VSS.t33 VSS.n311 272.676
R835 VSS.n145 VSS.n62 195
R836 VSS.n146 VSS.n145 195
R837 VSS.n160 VSS.n159 195
R838 VSS.n161 VSS.n160 195
R839 VSS.n58 VSS.n57 195
R840 VSS.n162 VSS.n58 195
R841 VSS.n59 VSS.n55 195
R842 VSS.n59 VSS.n53 195
R843 VSS.n182 VSS.n178 195
R844 VSS.n183 VSS.n182 195
R845 VSS.n186 VSS.n185 195
R846 VSS.n185 VSS.n184 195
R847 VSS.n48 VSS.n47 195
R848 VSS.n50 VSS.n48 195
R849 VSS.n49 VSS.n45 195
R850 VSS.n217 VSS.n49 195
R851 VSS.n231 VSS.n32 195
R852 VSS.n232 VSS.n231 195
R853 VSS.n246 VSS.n245 195
R854 VSS.n247 VSS.n246 195
R855 VSS.n28 VSS.n27 195
R856 VSS.n248 VSS.n28 195
R857 VSS.n29 VSS.n25 195
R858 VSS.n29 VSS.n23 195
R859 VSS.n268 VSS.n264 195
R860 VSS.n269 VSS.n268 195
R861 VSS.n284 VSS.n283 195
R862 VSS.n283 VSS.n282 195
R863 VSS.n280 VSS.n279 195
R864 VSS.n281 VSS.n280 195
R865 VSS.n274 VSS.n273 195
R866 VSS.n273 VSS.n272 195
R867 VSS.n98 VSS.n94 195
R868 VSS.n100 VSS.n98 195
R869 VSS.n99 VSS.n97 195
R870 VSS.n101 VSS.n99 195
R871 VSS.n78 VSS.n77 195
R872 VSS.n80 VSS.n78 195
R873 VSS.n79 VSS.n75 195
R874 VSS.n131 VSS.n79 195
R875 VSS.n314 VSS.n11 195
R876 VSS.n315 VSS.n314 195
R877 VSS.n330 VSS.n329 195
R878 VSS.n329 VSS.n328 195
R879 VSS.n326 VSS.n325 195
R880 VSS.n327 VSS.n326 195
R881 VSS.n320 VSS.n319 195
R882 VSS.n319 VSS.n318 195
R883 VSS VSS.n83 161.595
R884 VSS.n158 VSS.n60 146.25
R885 VSS.n60 VSS.t31 146.25
R886 VSS.n164 VSS.n163 146.25
R887 VSS.n163 VSS.t64 146.25
R888 VSS.n187 VSS.n180 146.25
R889 VSS.t17 VSS.n180 146.25
R890 VSS.n219 VSS.n218 146.25
R891 VSS.n218 VSS.t43 146.25
R892 VSS.n244 VSS.n30 146.25
R893 VSS.n30 VSS.t0 146.25
R894 VSS.n250 VSS.n249 146.25
R895 VSS.n249 VSS.t86 146.25
R896 VSS.n285 VSS.n266 146.25
R897 VSS.t93 VSS.n266 146.25
R898 VSS.n271 VSS.n270 146.25
R899 VSS.n270 VSS.t25 146.25
R900 VSS.n103 VSS.n102 146.25
R901 VSS.n102 VSS.t2 146.25
R902 VSS.n133 VSS.n132 146.25
R903 VSS.n132 VSS.t74 146.25
R904 VSS.n123 VSS.n122 146.25
R905 VSS.n124 VSS.n123 146.25
R906 VSS.n120 VSS.n89 146.25
R907 VSS.n111 VSS.n89 146.25
R908 VSS.n108 VSS.n90 146.25
R909 VSS.n112 VSS.n108 146.25
R910 VSS.n109 VSS.n107 146.25
R911 VSS.n113 VSS.n109 146.25
R912 VSS.n128 VSS.n74 146.25
R913 VSS.n129 VSS.n128 146.25
R914 VSS.n142 VSS.n141 146.25
R915 VSS.n143 VSS.n142 146.25
R916 VSS.n68 VSS.n67 146.25
R917 VSS.n144 VSS.n68 146.25
R918 VSS.n69 VSS.n63 146.25
R919 VSS.n148 VSS.n69 146.25
R920 VSS.n207 VSS.n206 146.25
R921 VSS.n208 VSS.n207 146.25
R922 VSS.n204 VSS.n173 146.25
R923 VSS.n195 VSS.n173 146.25
R924 VSS.n192 VSS.n174 146.25
R925 VSS.n196 VSS.n192 146.25
R926 VSS.n193 VSS.n191 146.25
R927 VSS.n197 VSS.n193 146.25
R928 VSS.n214 VSS.n44 146.25
R929 VSS.n215 VSS.n214 146.25
R930 VSS.n228 VSS.n227 146.25
R931 VSS.n229 VSS.n228 146.25
R932 VSS.n38 VSS.n37 146.25
R933 VSS.n230 VSS.n38 146.25
R934 VSS.n39 VSS.n33 146.25
R935 VSS.n234 VSS.n39 146.25
R936 VSS.n305 VSS.n304 146.25
R937 VSS.n306 VSS.n305 146.25
R938 VSS.n302 VSS.n259 146.25
R939 VSS.n293 VSS.n259 146.25
R940 VSS.n290 VSS.n260 146.25
R941 VSS.n294 VSS.n290 146.25
R942 VSS.n291 VSS.n289 146.25
R943 VSS.n295 VSS.n291 146.25
R944 VSS.n331 VSS.n13 146.25
R945 VSS.t105 VSS.n13 146.25
R946 VSS.n324 VSS.n15 146.25
R947 VSS.n15 VSS.t103 146.25
R948 VSS.n18 VSS.n4 146.25
R949 VSS.n19 VSS.n18 146.25
R950 VSS.n343 VSS.n342 146.25
R951 VSS.n342 VSS.n341 146.25
R952 VSS.n339 VSS.n338 146.25
R953 VSS.n340 VSS.n339 146.25
R954 VSS.n312 VSS.n10 146.25
R955 VSS.n313 VSS.n312 146.25
R956 VSS.n344 VSS.n343 105.695
R957 VSS.n344 VSS.n4 105.695
R958 VSS.n74 VSS.n71 105.695
R959 VSS.n141 VSS.n71 105.695
R960 VSS.n151 VSS.n67 105.695
R961 VSS.n151 VSS.n63 105.695
R962 VSS.n206 VSS.n205 105.695
R963 VSS.n205 VSS.n204 105.695
R964 VSS.n200 VSS.n174 105.695
R965 VSS.n200 VSS.n191 105.695
R966 VSS.n44 VSS.n41 105.695
R967 VSS.n227 VSS.n41 105.695
R968 VSS.n237 VSS.n37 105.695
R969 VSS.n237 VSS.n33 105.695
R970 VSS.n304 VSS.n303 105.695
R971 VSS.n303 VSS.n302 105.695
R972 VSS.n298 VSS.n260 105.695
R973 VSS.n298 VSS.n289 105.695
R974 VSS.n122 VSS.n121 105.695
R975 VSS.n121 VSS.n120 105.695
R976 VSS.n116 VSS.n90 105.695
R977 VSS.n116 VSS.n107 105.695
R978 VSS.n338 VSS.n7 105.695
R979 VSS.n10 VSS.n7 105.695
R980 VSS.n12 VSS.t106 84.1574
R981 VSS.n322 VSS.t104 84.1574
R982 VSS.n95 VSS.t3 84.1574
R983 VSS.n135 VSS.t75 84.1574
R984 VSS.n156 VSS.t32 84.1574
R985 VSS.n166 VSS.t65 84.1574
R986 VSS.n179 VSS.t18 84.1574
R987 VSS.n221 VSS.t44 84.1574
R988 VSS.n242 VSS.t1 84.1574
R989 VSS.n252 VSS.t87 84.1574
R990 VSS.n265 VSS.t94 84.1574
R991 VSS.n276 VSS.t26 84.1574
R992 VSS.n2 VSS.t50 83.7172
R993 VSS.n9 VSS.t10 83.7172
R994 VSS.n73 VSS.t99 83.7172
R995 VSS.n65 VSS.t20 83.7172
R996 VSS.n170 VSS.t40 83.7172
R997 VSS.n176 VSS.t42 83.7172
R998 VSS.n43 VSS.t69 83.7172
R999 VSS.n35 VSS.t5 83.7172
R1000 VSS.n256 VSS.t36 83.7172
R1001 VSS.n262 VSS.t28 83.7172
R1002 VSS.n86 VSS.t83 83.7172
R1003 VSS.n92 VSS.t73 83.7172
R1004 VSS.n2 VSS.n1 75.905
R1005 VSS.n9 VSS.n8 75.905
R1006 VSS.n73 VSS.n72 75.905
R1007 VSS.n65 VSS.n64 75.905
R1008 VSS.n170 VSS.n169 75.905
R1009 VSS.n176 VSS.n175 75.905
R1010 VSS.n43 VSS.n42 75.905
R1011 VSS.n35 VSS.n34 75.905
R1012 VSS.n256 VSS.n255 75.905
R1013 VSS.n262 VSS.n261 75.905
R1014 VSS.n86 VSS.n85 75.905
R1015 VSS.n92 VSS.n91 75.905
R1016 VSS.n121 VSS.n82 73.1255
R1017 VSS.n110 VSS.n82 73.1255
R1018 VSS.n116 VSS.n115 73.1255
R1019 VSS.n115 VSS.n114 73.1255
R1020 VSS.n71 VSS.n70 73.1255
R1021 VSS.n127 VSS.n70 73.1255
R1022 VSS.n151 VSS.n150 73.1255
R1023 VSS.n150 VSS.n149 73.1255
R1024 VSS.n205 VSS.n54 73.1255
R1025 VSS.n194 VSS.n54 73.1255
R1026 VSS.n200 VSS.n199 73.1255
R1027 VSS.n199 VSS.n198 73.1255
R1028 VSS.n41 VSS.n40 73.1255
R1029 VSS.n213 VSS.n40 73.1255
R1030 VSS.n237 VSS.n236 73.1255
R1031 VSS.n236 VSS.n235 73.1255
R1032 VSS.n303 VSS.n24 73.1255
R1033 VSS.n292 VSS.n24 73.1255
R1034 VSS.n298 VSS.n297 73.1255
R1035 VSS.n297 VSS.n296 73.1255
R1036 VSS.n344 VSS.n5 73.1255
R1037 VSS.n17 VSS.n5 73.1255
R1038 VSS.n7 VSS.n6 73.1255
R1039 VSS.n311 VSS.n6 73.1255
R1040 VSS.n133 VSS.n77 68.7561
R1041 VSS.n133 VSS.n75 68.7561
R1042 VSS.n159 VSS.n158 68.7561
R1043 VSS.n158 VSS.n62 68.7561
R1044 VSS.n164 VSS.n57 68.7561
R1045 VSS.n164 VSS.n55 68.7561
R1046 VSS.n187 VSS.n186 68.7561
R1047 VSS.n187 VSS.n178 68.7561
R1048 VSS.n219 VSS.n47 68.7561
R1049 VSS.n219 VSS.n45 68.7561
R1050 VSS.n245 VSS.n244 68.7561
R1051 VSS.n244 VSS.n32 68.7561
R1052 VSS.n250 VSS.n27 68.7561
R1053 VSS.n250 VSS.n25 68.7561
R1054 VSS.n285 VSS.n284 68.7561
R1055 VSS.n285 VSS.n264 68.7561
R1056 VSS.n279 VSS.n271 68.7561
R1057 VSS.n274 VSS.n271 68.7561
R1058 VSS.n103 VSS.n97 68.7561
R1059 VSS.n103 VSS.n94 68.7561
R1060 VSS.n324 VSS.n320 68.7561
R1061 VSS.n325 VSS.n324 68.7561
R1062 VSS.n331 VSS.n330 68.7561
R1063 VSS.n331 VSS.n11 68.7561
R1064 VSS.n1 VSS.t63 17.4005
R1065 VSS.n1 VSS.t97 17.4005
R1066 VSS.n8 VSS.t108 17.4005
R1067 VSS.n8 VSS.t34 17.4005
R1068 VSS.n72 VSS.t57 17.4005
R1069 VSS.n72 VSS.t89 17.4005
R1070 VSS.n64 VSS.t12 17.4005
R1071 VSS.n64 VSS.t53 17.4005
R1072 VSS.n169 VSS.t59 17.4005
R1073 VSS.n169 VSS.t91 17.4005
R1074 VSS.n175 VSS.t38 17.4005
R1075 VSS.n175 VSS.t55 17.4005
R1076 VSS.n42 VSS.t67 17.4005
R1077 VSS.n42 VSS.t71 17.4005
R1078 VSS.n34 VSS.t22 17.4005
R1079 VSS.n34 VSS.t7 17.4005
R1080 VSS.n255 VSS.t46 17.4005
R1081 VSS.n255 VSS.t48 17.4005
R1082 VSS.n261 VSS.t24 17.4005
R1083 VSS.n261 VSS.t30 17.4005
R1084 VSS.n85 VSS.t81 17.4005
R1085 VSS.n85 VSS.t85 17.4005
R1086 VSS.n91 VSS.t79 17.4005
R1087 VSS.n91 VSS.t77 17.4005
R1088 VSS.n105 VSS.n94 3.46248
R1089 VSS.n77 VSS.n76 3.46248
R1090 VSS.n136 VSS.n75 3.46248
R1091 VSS.n57 VSS.n56 3.46248
R1092 VSS.n155 VSS.n62 3.46248
R1093 VSS.n159 VSS.n61 3.46248
R1094 VSS.n167 VSS.n55 3.46248
R1095 VSS.n47 VSS.n46 3.46248
R1096 VSS.n189 VSS.n178 3.46248
R1097 VSS.n186 VSS.n181 3.46248
R1098 VSS.n222 VSS.n45 3.46248
R1099 VSS.n27 VSS.n26 3.46248
R1100 VSS.n241 VSS.n32 3.46248
R1101 VSS.n245 VSS.n31 3.46248
R1102 VSS.n253 VSS.n25 3.46248
R1103 VSS.n279 VSS.n278 3.46248
R1104 VSS.n287 VSS.n264 3.46248
R1105 VSS.n284 VSS.n267 3.46248
R1106 VSS.n275 VSS.n274 3.46248
R1107 VSS.n97 VSS.n96 3.46248
R1108 VSS.n325 VSS.n16 3.46248
R1109 VSS.n321 VSS.n320 3.46248
R1110 VSS.n333 VSS.n11 3.46248
R1111 VSS.n330 VSS.n14 3.46248
R1112 VSS.n338 VSS.n337 2.82278
R1113 VSS.n4 VSS.n0 2.82278
R1114 VSS.n343 VSS.n3 2.82278
R1115 VSS.n137 VSS.n74 2.82278
R1116 VSS.n141 VSS.n140 2.82278
R1117 VSS.n67 VSS.n66 2.82278
R1118 VSS.n154 VSS.n63 2.82278
R1119 VSS.n206 VSS.n168 2.82278
R1120 VSS.n204 VSS.n203 2.82278
R1121 VSS.n202 VSS.n174 2.82278
R1122 VSS.n191 VSS.n190 2.82278
R1123 VSS.n223 VSS.n44 2.82278
R1124 VSS.n227 VSS.n226 2.82278
R1125 VSS.n37 VSS.n36 2.82278
R1126 VSS.n240 VSS.n33 2.82278
R1127 VSS.n304 VSS.n254 2.82278
R1128 VSS.n302 VSS.n301 2.82278
R1129 VSS.n300 VSS.n260 2.82278
R1130 VSS.n289 VSS.n288 2.82278
R1131 VSS.n122 VSS.n84 2.82278
R1132 VSS.n120 VSS.n119 2.82278
R1133 VSS.n118 VSS.n90 2.82278
R1134 VSS.n107 VSS.n106 2.82278
R1135 VSS.n334 VSS.n10 2.82278
R1136 VSS.n286 VSS.n285 2.3255
R1137 VSS.n277 VSS.n271 2.3255
R1138 VSS.n244 VSS.n243 2.3255
R1139 VSS.n251 VSS.n250 2.3255
R1140 VSS.n188 VSS.n187 2.3255
R1141 VSS.n220 VSS.n219 2.3255
R1142 VSS.n158 VSS.n157 2.3255
R1143 VSS.n165 VSS.n164 2.3255
R1144 VSS.n134 VSS.n133 2.3255
R1145 VSS.n104 VSS.n103 2.3255
R1146 VSS.n332 VSS.n331 2.3255
R1147 VSS.n324 VSS.n323 2.3255
R1148 VSS.n303 VSS.n258 1.32907
R1149 VSS.n299 VSS.n298 1.32907
R1150 VSS.n225 VSS.n41 1.32907
R1151 VSS.n238 VSS.n237 1.32907
R1152 VSS.n205 VSS.n172 1.32907
R1153 VSS.n201 VSS.n200 1.32907
R1154 VSS.n139 VSS.n71 1.32907
R1155 VSS.n152 VSS.n151 1.32907
R1156 VSS.n121 VSS.n88 1.32907
R1157 VSS.n117 VSS.n116 1.32907
R1158 VSS.n345 VSS.n344 1.32907
R1159 VSS.n336 VSS.n7 1.32907
R1160 VSS.n84 VSS 0.90794
R1161 VSS.n346 VSS.n2 0.685283
R1162 VSS.n335 VSS.n9 0.685283
R1163 VSS.n138 VSS.n73 0.685283
R1164 VSS.n153 VSS.n65 0.685283
R1165 VSS.n171 VSS.n170 0.685283
R1166 VSS.n177 VSS.n176 0.685283
R1167 VSS.n224 VSS.n43 0.685283
R1168 VSS.n239 VSS.n35 0.685283
R1169 VSS.n257 VSS.n256 0.685283
R1170 VSS.n263 VSS.n262 0.685283
R1171 VSS.n87 VSS.n86 0.685283
R1172 VSS.n93 VSS.n92 0.685283
R1173 VSS.n275 VSS 0.479667
R1174 VSS VSS.n253 0.479667
R1175 VSS VSS.n222 0.479667
R1176 VSS VSS.n167 0.479667
R1177 VSS VSS.n136 0.479667
R1178 VSS VSS.n287 0.466646
R1179 VSS.n241 VSS 0.466646
R1180 VSS VSS.n189 0.466646
R1181 VSS.n155 VSS 0.466646
R1182 VSS VSS.n105 0.466646
R1183 VSS VSS.n333 0.466646
R1184 VSS.n301 VSS.n300 0.430188
R1185 VSS.n226 VSS.n36 0.430188
R1186 VSS.n203 VSS.n202 0.430188
R1187 VSS.n140 VSS.n66 0.430188
R1188 VSS.n119 VSS.n118 0.430188
R1189 VSS.n337 VSS.n3 0.430188
R1190 VSS.n321 VSS 0.404146
R1191 VSS.n301 VSS.n258 0.359875
R1192 VSS.n300 VSS.n299 0.359875
R1193 VSS.n226 VSS.n225 0.359875
R1194 VSS.n238 VSS.n36 0.359875
R1195 VSS.n203 VSS.n172 0.359875
R1196 VSS.n202 VSS.n201 0.359875
R1197 VSS.n140 VSS.n139 0.359875
R1198 VSS.n152 VSS.n66 0.359875
R1199 VSS.n119 VSS.n88 0.359875
R1200 VSS.n118 VSS.n117 0.359875
R1201 VSS.n345 VSS.n3 0.359875
R1202 VSS.n337 VSS.n336 0.359875
R1203 VSS.n258 VSS.n257 0.229667
R1204 VSS.n299 VSS.n263 0.229667
R1205 VSS.n225 VSS.n224 0.229667
R1206 VSS.n239 VSS.n238 0.229667
R1207 VSS.n172 VSS.n171 0.229667
R1208 VSS.n201 VSS.n177 0.229667
R1209 VSS.n139 VSS.n138 0.229667
R1210 VSS.n153 VSS.n152 0.229667
R1211 VSS.n88 VSS.n87 0.229667
R1212 VSS.n117 VSS.n93 0.229667
R1213 VSS.n346 VSS.n345 0.229667
R1214 VSS.n336 VSS.n335 0.229667
R1215 VSS.n254 VSS 0.191906
R1216 VSS.n223 VSS 0.191906
R1217 VSS.n168 VSS 0.191906
R1218 VSS.n137 VSS 0.191906
R1219 VSS VSS.n0 0.191906
R1220 VSS.n287 VSS.n286 0.189302
R1221 VSS.n278 VSS.n277 0.189302
R1222 VSS.n243 VSS.n241 0.189302
R1223 VSS.n251 VSS.n26 0.189302
R1224 VSS.n189 VSS.n188 0.189302
R1225 VSS.n220 VSS.n46 0.189302
R1226 VSS.n157 VSS.n155 0.189302
R1227 VSS.n165 VSS.n56 0.189302
R1228 VSS.n105 VSS.n104 0.189302
R1229 VSS.n134 VSS.n76 0.189302
R1230 VSS.n333 VSS.n332 0.189302
R1231 VSS.n323 VSS.n16 0.189302
R1232 VSS.n278 VSS.n267 0.141125
R1233 VSS.n31 VSS.n26 0.141125
R1234 VSS.n181 VSS.n46 0.141125
R1235 VSS.n61 VSS.n56 0.141125
R1236 VSS.n96 VSS.n76 0.141125
R1237 VSS.n16 VSS.n14 0.141125
R1238 VSS.n267 VSS.n265 0.13201
R1239 VSS.n276 VSS.n275 0.13201
R1240 VSS.n242 VSS.n31 0.13201
R1241 VSS.n253 VSS.n252 0.13201
R1242 VSS.n181 VSS.n179 0.13201
R1243 VSS.n222 VSS.n221 0.13201
R1244 VSS.n156 VSS.n61 0.13201
R1245 VSS.n167 VSS.n166 0.13201
R1246 VSS.n96 VSS.n95 0.13201
R1247 VSS.n136 VSS.n135 0.13201
R1248 VSS.n14 VSS.n12 0.13201
R1249 VSS.n322 VSS.n321 0.13201
R1250 VSS.n288 VSS.n263 0.130708
R1251 VSS.n240 VSS.n239 0.130708
R1252 VSS.n190 VSS.n177 0.130708
R1253 VSS.n154 VSS.n153 0.130708
R1254 VSS.n106 VSS.n93 0.130708
R1255 VSS.n335 VSS.n334 0.130708
R1256 VSS.n257 VSS 0.124198
R1257 VSS.n224 VSS 0.124198
R1258 VSS.n171 VSS 0.124198
R1259 VSS.n138 VSS 0.124198
R1260 VSS.n87 VSS 0.124198
R1261 VSS VSS.n346 0.124198
R1262 VSS.n288 VSS 0.0695104
R1263 VSS VSS.n240 0.0695104
R1264 VSS.n190 VSS 0.0695104
R1265 VSS VSS.n154 0.0695104
R1266 VSS.n106 VSS 0.0695104
R1267 VSS.n334 VSS 0.0695104
R1268 VSS.n286 VSS.n265 0.0577917
R1269 VSS.n277 VSS.n276 0.0577917
R1270 VSS.n243 VSS.n242 0.0577917
R1271 VSS.n252 VSS.n251 0.0577917
R1272 VSS.n188 VSS.n179 0.0577917
R1273 VSS.n221 VSS.n220 0.0577917
R1274 VSS.n157 VSS.n156 0.0577917
R1275 VSS.n166 VSS.n165 0.0577917
R1276 VSS.n104 VSS.n95 0.0577917
R1277 VSS.n135 VSS.n134 0.0577917
R1278 VSS.n332 VSS.n12 0.0577917
R1279 VSS.n323 VSS.n322 0.0577917
R1280 VSS VSS.n254 0.00701042
R1281 VSS VSS.n223 0.00701042
R1282 VSS VSS.n168 0.00701042
R1283 VSS VSS.n137 0.00701042
R1284 VSS VSS.n84 0.00701042
R1285 VSS VSS.n0 0.00701042
R1286 variable_delay_unit_3.in.n0 variable_delay_unit_3.in.t4 607.409
R1287 variable_delay_unit_3.in.n2 variable_delay_unit_3.in.t2 543.053
R1288 variable_delay_unit_3.in.n0 variable_delay_unit_3.in.t5 321.423
R1289 variable_delay_unit_3.in variable_delay_unit_3.in.n2 221.778
R1290 variable_delay_unit_3.in.n2 variable_delay_unit_3.in.t3 221.72
R1291 variable_delay_unit_3.in variable_delay_unit_3.in.n0 161.72
R1292 variable_delay_unit_3.in.n1 variable_delay_unit_3.in.t1 84.7227
R1293 variable_delay_unit_3.in.n1 variable_delay_unit_3.in.t0 84.0867
R1294 variable_delay_unit_3.in.n3 variable_delay_unit_3.in 20.0791
R1295 variable_delay_unit_3.in variable_delay_unit_3.in.n3 0.851271
R1296 variable_delay_unit_3.in.n3 variable_delay_unit_3.in.n1 0.465495
R1297 variable_delay_unit_4.in.n0 variable_delay_unit_4.in.t3 607.409
R1298 variable_delay_unit_4.in.n2 variable_delay_unit_4.in.t2 543.053
R1299 variable_delay_unit_4.in.n0 variable_delay_unit_4.in.t5 321.423
R1300 variable_delay_unit_4.in variable_delay_unit_4.in.n2 221.778
R1301 variable_delay_unit_4.in.n2 variable_delay_unit_4.in.t4 221.72
R1302 variable_delay_unit_4.in variable_delay_unit_4.in.n0 161.72
R1303 variable_delay_unit_4.in.n1 variable_delay_unit_4.in.t1 84.7227
R1304 variable_delay_unit_4.in.n1 variable_delay_unit_4.in.t0 84.0867
R1305 variable_delay_unit_4.in.n3 variable_delay_unit_4.in 20.0791
R1306 variable_delay_unit_4.in variable_delay_unit_4.in.n3 0.851271
R1307 variable_delay_unit_4.in.n3 variable_delay_unit_4.in.n1 0.465495
R1308 variable_delay_unit_2.in.n0 variable_delay_unit_2.in.t4 607.409
R1309 variable_delay_unit_2.in.n2 variable_delay_unit_2.in.t2 543.053
R1310 variable_delay_unit_2.in.n0 variable_delay_unit_2.in.t5 321.423
R1311 variable_delay_unit_2.in variable_delay_unit_2.in.n2 221.778
R1312 variable_delay_unit_2.in.n2 variable_delay_unit_2.in.t3 221.72
R1313 variable_delay_unit_2.in variable_delay_unit_2.in.n0 161.72
R1314 variable_delay_unit_2.in.n1 variable_delay_unit_2.in.t0 84.7227
R1315 variable_delay_unit_2.in.n1 variable_delay_unit_2.in.t1 84.0867
R1316 variable_delay_unit_2.in.n3 variable_delay_unit_2.in 20.0791
R1317 variable_delay_unit_2.in variable_delay_unit_2.in.n3 0.851271
R1318 variable_delay_unit_2.in.n3 variable_delay_unit_2.in.n1 0.465495
R1319 en_0.n2 en_0.t0 628.097
R1320 en_0.n3 en_0.t6 622.766
R1321 en_0.n0 en_0.t1 543.053
R1322 en_0.n2 en_0.t4 523.774
R1323 en_0.n1 en_0.t3 304.647
R1324 en_0.n1 en_0.t5 304.647
R1325 en_0.n0 en_0.t2 221.72
R1326 en_0.n5 en_0.n0 220.263
R1327 en_0.n1 en_0.t7 202.44
R1328 en_0 en_0.n1 168.969
R1329 en_0 en_0.n3 166.147
R1330 en_0 en_0.n4 3.17729
R1331 en_0.n4 en_0 1.40175
R1332 en_0.n3 en_0.n2 1.09595
R1333 en_0.n4 en_0 0.443357
R1334 en_0.n5 en_0 0.088
R1335 en_0 en_0.n5 0.063
R1336 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t6 628.097
R1337 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.t7 622.766
R1338 variable_delay_unit_1.tristate_inverter_1.en.n3 variable_delay_unit_1.tristate_inverter_1.en.t4 523.774
R1339 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t3 304.647
R1340 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t2 304.647
R1341 variable_delay_unit_1.tristate_inverter_1.en.n0 variable_delay_unit_1.tristate_inverter_1.en.t5 202.44
R1342 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n0 168.969
R1343 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n4 166.147
R1344 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t1 84.7557
R1345 variable_delay_unit_1.tristate_inverter_1.en.n1 variable_delay_unit_1.tristate_inverter_1.en.t0 84.1197
R1346 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en.n1 12.6535
R1347 variable_delay_unit_1.tristate_inverter_1.en.n2 variable_delay_unit_1.tristate_inverter_1.en 5.58443
R1348 variable_delay_unit_1.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en.n2 4.59003
R1349 variable_delay_unit_1.tristate_inverter_1.en.n4 variable_delay_unit_1.tristate_inverter_1.en.n3 1.09595
R1350 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t3 628.097
R1351 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.t5 622.766
R1352 variable_delay_unit_0.tristate_inverter_1.en.n3 variable_delay_unit_0.tristate_inverter_1.en.t7 523.774
R1353 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t6 304.647
R1354 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t2 304.647
R1355 variable_delay_unit_0.tristate_inverter_1.en.n0 variable_delay_unit_0.tristate_inverter_1.en.t4 202.44
R1356 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n0 168.969
R1357 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n4 166.147
R1358 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t1 84.7557
R1359 variable_delay_unit_0.tristate_inverter_1.en.n1 variable_delay_unit_0.tristate_inverter_1.en.t0 84.1197
R1360 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en.n1 12.6535
R1361 variable_delay_unit_0.tristate_inverter_1.en.n2 variable_delay_unit_0.tristate_inverter_1.en 5.58443
R1362 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_0.tristate_inverter_1.en.n2 4.59003
R1363 variable_delay_unit_0.tristate_inverter_1.en.n4 variable_delay_unit_0.tristate_inverter_1.en.n3 1.09595
R1364 variable_delay_unit_5.in.n0 variable_delay_unit_5.in.t4 607.409
R1365 variable_delay_unit_5.in.n2 variable_delay_unit_5.in.t2 543.053
R1366 variable_delay_unit_5.in.n0 variable_delay_unit_5.in.t5 321.423
R1367 variable_delay_unit_5.in variable_delay_unit_5.in.n2 221.778
R1368 variable_delay_unit_5.in.n2 variable_delay_unit_5.in.t3 221.72
R1369 variable_delay_unit_5.in variable_delay_unit_5.in.n0 161.72
R1370 variable_delay_unit_5.in.n1 variable_delay_unit_5.in.t1 84.7227
R1371 variable_delay_unit_5.in.n1 variable_delay_unit_5.in.t0 84.0867
R1372 variable_delay_unit_5.in.n3 variable_delay_unit_5.in 20.0791
R1373 variable_delay_unit_5.in variable_delay_unit_5.in.n3 0.851271
R1374 variable_delay_unit_5.in.n3 variable_delay_unit_5.in.n1 0.465495
R1375 variable_delay_unit_5.forward.n0 variable_delay_unit_5.forward.t2 607.409
R1376 variable_delay_unit_5.forward.n0 variable_delay_unit_5.forward.t3 321.423
R1377 variable_delay_unit_5.forward variable_delay_unit_5.forward.n0 161.72
R1378 variable_delay_unit_5.forward.n1 variable_delay_unit_5.forward.t1 84.7227
R1379 variable_delay_unit_5.forward.n1 variable_delay_unit_5.forward.t0 84.0867
R1380 variable_delay_unit_5.forward.n2 variable_delay_unit_5.forward 19.8934
R1381 variable_delay_unit_5.forward variable_delay_unit_5.forward.n2 0.851271
R1382 variable_delay_unit_5.forward.n2 variable_delay_unit_5.forward.n1 0.465495
R1383 en_4.n0 en_4.t2 628.097
R1384 en_4.n1 en_4.t0 622.766
R1385 en_4.n2 en_4.t5 543.053
R1386 en_4.n0 en_4.t4 523.774
R1387 en_4.n4 en_4.t3 304.647
R1388 en_4.n4 en_4.t7 304.647
R1389 en_4.n2 en_4.t6 221.72
R1390 en_4 en_4.n2 220.304
R1391 en_4.n4 en_4.t1 202.44
R1392 en_4 en_4.n4 168.969
R1393 en_4 en_4.n1 166.147
R1394 en_4.n3 en_4 3.22371
R1395 en_4.n3 en_4 1.40175
R1396 en_4.n1 en_4.n0 1.09595
R1397 en_4 en_4.n3 0.443357
R1398 en_3.n2 en_3.t0 628.097
R1399 en_3.n3 en_3.t7 622.766
R1400 en_3.n0 en_3.t3 543.053
R1401 en_3.n2 en_3.t2 523.774
R1402 en_3.n1 en_3.t5 304.647
R1403 en_3.n1 en_3.t6 304.647
R1404 en_3.n0 en_3.t4 221.72
R1405 en_3.n5 en_3.n0 220.263
R1406 en_3.n1 en_3.t1 202.44
R1407 en_3 en_3.n1 168.969
R1408 en_3 en_3.n3 166.147
R1409 en_3 en_3.n4 3.15229
R1410 en_3.n4 en_3 1.40175
R1411 en_3.n3 en_3.n2 1.09595
R1412 en_3.n4 en_3 0.443357
R1413 en_3.n5 en_3 0.113
R1414 en_3 en_3.n5 0.063
R1415 en_2.n2 en_2.t1 628.097
R1416 en_2.n3 en_2.t7 622.766
R1417 en_2.n0 en_2.t3 543.053
R1418 en_2.n2 en_2.t4 523.774
R1419 en_2.n1 en_2.t2 304.647
R1420 en_2.n1 en_2.t6 304.647
R1421 en_2.n0 en_2.t5 221.72
R1422 en_2.n5 en_2.n0 220.263
R1423 en_2.n1 en_2.t0 202.44
R1424 en_2 en_2.n1 168.969
R1425 en_2 en_2.n3 166.147
R1426 en_2 en_2.n4 3.09157
R1427 en_2.n4 en_2 1.40175
R1428 en_2.n3 en_2.n2 1.09595
R1429 en_2.n4 en_2 0.443357
R1430 en_2.n5 en_2 0.173714
R1431 en_2 en_2.n5 0.063
R1432 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t2 607.409
R1433 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t4 543.053
R1434 variable_delay_unit_1.in.n0 variable_delay_unit_1.in.t3 321.423
R1435 variable_delay_unit_1.in variable_delay_unit_1.in.n2 221.778
R1436 variable_delay_unit_1.in.n2 variable_delay_unit_1.in.t5 221.72
R1437 variable_delay_unit_1.in variable_delay_unit_1.in.n0 161.72
R1438 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t0 84.7227
R1439 variable_delay_unit_1.in.n1 variable_delay_unit_1.in.t1 84.0867
R1440 variable_delay_unit_1.in.n3 variable_delay_unit_1.in 20.0791
R1441 variable_delay_unit_1.in variable_delay_unit_1.in.n3 0.851271
R1442 variable_delay_unit_1.in.n3 variable_delay_unit_1.in.n1 0.465495
R1443 out.n0 out.t1 84.8477
R1444 out.n2 out.t2 84.8477
R1445 out.n0 out.t0 84.2063
R1446 out.n2 out.t3 84.1683
R1447 out out.n3 10.0241
R1448 out.n1 out 0.681535
R1449 out out.n0 0.287138
R1450 out.n3 out 0.0803611
R1451 out.n3 out.n2 0.0508472
R1452 out.n1 out 0.013431
R1453 out out.n1 0.0109167
R1454 variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_unit_4.tristate_inverter_1.en.t5 628.097
R1455 variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_unit_4.tristate_inverter_1.en.t7 622.766
R1456 variable_delay_unit_4.tristate_inverter_1.en.n3 variable_delay_unit_4.tristate_inverter_1.en.t3 523.774
R1457 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t2 304.647
R1458 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t4 304.647
R1459 variable_delay_unit_4.tristate_inverter_1.en.n0 variable_delay_unit_4.tristate_inverter_1.en.t6 202.44
R1460 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n0 168.969
R1461 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n4 166.147
R1462 variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_unit_4.tristate_inverter_1.en.t1 84.7557
R1463 variable_delay_unit_4.tristate_inverter_1.en.n1 variable_delay_unit_4.tristate_inverter_1.en.t0 84.1197
R1464 variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_unit_4.tristate_inverter_1.en.n1 12.6535
R1465 variable_delay_unit_4.tristate_inverter_1.en.n2 variable_delay_unit_4.tristate_inverter_1.en 5.58443
R1466 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en.n2 4.59003
R1467 variable_delay_unit_4.tristate_inverter_1.en.n4 variable_delay_unit_4.tristate_inverter_1.en.n3 1.09595
R1468 variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_unit_3.tristate_inverter_1.en.t5 628.097
R1469 variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_unit_3.tristate_inverter_1.en.t6 622.766
R1470 variable_delay_unit_3.tristate_inverter_1.en.n3 variable_delay_unit_3.tristate_inverter_1.en.t3 523.774
R1471 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t7 304.647
R1472 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t2 304.647
R1473 variable_delay_unit_3.tristate_inverter_1.en.n0 variable_delay_unit_3.tristate_inverter_1.en.t4 202.44
R1474 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n0 168.969
R1475 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n4 166.147
R1476 variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_unit_3.tristate_inverter_1.en.t1 84.7557
R1477 variable_delay_unit_3.tristate_inverter_1.en.n1 variable_delay_unit_3.tristate_inverter_1.en.t0 84.1197
R1478 variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_unit_3.tristate_inverter_1.en.n1 12.6535
R1479 variable_delay_unit_3.tristate_inverter_1.en.n2 variable_delay_unit_3.tristate_inverter_1.en 5.58443
R1480 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_3.tristate_inverter_1.en.n2 4.59003
R1481 variable_delay_unit_3.tristate_inverter_1.en.n4 variable_delay_unit_3.tristate_inverter_1.en.n3 1.09595
R1482 in.n0 in.t0 543.053
R1483 in.n0 in.t1 221.72
R1484 in in.n0 221.565
C0 VDD variable_delay_unit_1.out 1.34424f
C1 a_14288_772# variable_delay_unit_4.out 0.493816f
C2 a_17236_352# variable_delay_unit_5.out 0.172055f
C3 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_5.out 0.085059f
C4 a_8392_352# en_2 0.001909f
C5 variable_delay_unit_3.tristate_inverter_1.en en_4 9.38e-20
C6 en_2 a_5444_772# 6.99e-20
C7 variable_delay_unit_3.in a_7510_352# 0.054206f
C8 en_2 en_3 0.010459f
C9 variable_delay_unit_2.in variable_delay_unit_2.out 0.499092f
C10 a_11340_772# variable_delay_unit_3.tristate_inverter_1.en 0.029284f
C11 variable_delay_unit_3.in en_2 0.574722f
C12 en_2 variable_delay_unit_4.in 3.37e-20
C13 a_16354_772# variable_delay_unit_5.forward 0.088132f
C14 en_2 en_1 0.010459f
C15 a_2496_352# en_0 0.001909f
C16 a_14288_772# variable_delay_unit_5.in 0.020173f
C17 VDD variable_delay_unit_2.in 2.12807f
C18 a_5444_352# variable_delay_unit_2.out 0.070146f
C19 in en_0 0.259572f
C20 en_2 variable_delay_unit_3.out 0.043504f
C21 variable_delay_unit_2.in variable_delay_unit_1.out 0.235667f
C22 a_2496_772# en_0 0.124274f
C23 variable_delay_unit_5.in variable_delay_unit_5.forward 0.087283f
C24 en_3 variable_delay_unit_4.tristate_inverter_1.en 1.5e-19
C25 variable_delay_unit_4.out variable_delay_unit_5.tristate_inverter_1.en 0.002141f
C26 VDD a_5444_352# 0.001468f
C27 variable_delay_unit_4.in variable_delay_unit_4.tristate_inverter_1.en 0.09141f
C28 en_0 variable_delay_unit_1.tristate_inverter_1.en 1.5e-19
C29 VDD a_4562_772# 1.6584f
C30 a_14288_772# a_14288_352# 0.011184f
C31 a_13406_772# variable_delay_unit_4.out 0.505512f
C32 a_16354_772# variable_delay_unit_5.tristate_inverter_1.en 0.11539f
C33 variable_delay_unit_2.out variable_delay_unit_2.tristate_inverter_1.en 0.12029f
C34 variable_delay_unit_3.in a_7510_772# 0.088132f
C35 a_5444_352# variable_delay_unit_1.out 0.172055f
C36 variable_delay_unit_4.out variable_delay_unit_5.out 0.071795f
C37 variable_delay_unit_1.out a_4562_772# 0.505512f
C38 variable_delay_unit_1.in variable_delay_unit_0.tristate_inverter_1.en 0.814958f
C39 out en_0 0.218964f
C40 a_16354_772# variable_delay_unit_5.out 0.505512f
C41 VDD a_2496_352# 0.001468f
C42 en_1 variable_delay_unit_0.tristate_inverter_1.en 9.38e-20
C43 VDD a_14288_772# 1.65847f
C44 variable_delay_unit_2.out variable_delay_unit_1.tristate_inverter_1.en 0.085059f
C45 en_2 variable_delay_unit_3.tristate_inverter_1.en 1.5e-19
C46 a_13406_352# variable_delay_unit_4.tristate_inverter_1.en 2.39e-19
C47 VDD in 0.238594f
C48 VDD variable_delay_unit_2.tristate_inverter_1.en 2.77611f
C49 a_2496_352# variable_delay_unit_1.out 0.070146f
C50 variable_delay_unit_3.out variable_delay_unit_4.tristate_inverter_1.en 0.002141f
C51 variable_delay_unit_1.in a_1614_772# 0.088132f
C52 variable_delay_unit_5.in variable_delay_unit_5.tristate_inverter_1.en 0.09141f
C53 variable_delay_unit_1.out variable_delay_unit_2.tristate_inverter_1.en 0.002141f
C54 variable_delay_unit_5.in a_13406_772# 0.088132f
C55 VDD a_2496_772# 1.6584f
C56 a_8392_772# variable_delay_unit_2.out 0.493816f
C57 a_1614_352# variable_delay_unit_0.tristate_inverter_1.en 2.39e-19
C58 VDD variable_delay_unit_5.forward 2.28561f
C59 variable_delay_unit_5.in variable_delay_unit_5.out 0.499092f
C60 variable_delay_unit_4.tristate_inverter_1.en en_4 1.09349f
C61 VDD variable_delay_unit_1.tristate_inverter_1.en 2.77611f
C62 variable_delay_unit_1.out a_2496_772# 0.071074f
C63 variable_delay_unit_2.in a_4562_772# 0.088132f
C64 variable_delay_unit_1.out variable_delay_unit_1.tristate_inverter_1.en 0.12029f
C65 a_1614_352# a_1614_772# 0.004142f
C66 en_3 a_10458_772# 0.042718f
C67 VDD out 1.15938f
C68 VDD a_8392_772# 1.6584f
C69 variable_delay_unit_3.in a_10458_772# 8.82e-20
C70 variable_delay_unit_4.in a_10458_772# 0.088132f
C71 a_17236_352# a_17236_772# 0.011184f
C72 en_3 variable_delay_unit_4.out 0.043504f
C73 variable_delay_unit_4.in variable_delay_unit_4.out 0.499092f
C74 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.tristate_inverter_1.en 0.002365f
C75 VDD a_4562_352# 6.98e-19
C76 variable_delay_unit_1.out out 0.071795f
C77 a_14288_352# variable_delay_unit_5.out 0.070146f
C78 variable_delay_unit_2.in variable_delay_unit_2.tristate_inverter_1.en 0.09141f
C79 en_3 a_11340_352# 0.001909f
C80 en_2 a_7510_352# 0.15982f
C81 a_16354_352# a_16354_772# 0.004142f
C82 variable_delay_unit_3.in a_11340_352# 7.65e-21
C83 variable_delay_unit_1.out a_4562_352# 0.222585f
C84 VDD variable_delay_unit_5.tristate_inverter_1.en 3.86957f
C85 VDD a_13406_772# 1.6584f
C86 variable_delay_unit_3.out a_10458_772# 0.505512f
C87 VDD variable_delay_unit_5.out 1.5668f
C88 a_13406_352# variable_delay_unit_4.out 0.222585f
C89 variable_delay_unit_2.in variable_delay_unit_1.tristate_inverter_1.en 0.814958f
C90 variable_delay_unit_3.out variable_delay_unit_4.out 0.071795f
C91 en_3 variable_delay_unit_5.in 3.37e-20
C92 variable_delay_unit_5.in variable_delay_unit_4.in 0.087283f
C93 a_16354_352# variable_delay_unit_5.in 8.82e-20
C94 variable_delay_unit_3.out a_11340_352# 0.172055f
C95 variable_delay_unit_2.in a_8392_772# 7.65e-21
C96 variable_delay_unit_4.out en_4 0.224474f
C97 variable_delay_unit_1.in en_0 0.574722f
C98 a_2496_352# in 7.65e-21
C99 en_3 a_10458_352# 0.15982f
C100 a_5444_352# variable_delay_unit_1.tristate_inverter_1.en 0.15982f
C101 variable_delay_unit_2.in a_4562_352# 0.054206f
C102 a_8392_352# variable_delay_unit_2.out 0.172055f
C103 variable_delay_unit_2.out a_5444_772# 0.071074f
C104 variable_delay_unit_3.in a_10458_352# 8.82e-20
C105 a_10458_352# variable_delay_unit_4.in 0.054206f
C106 a_4562_772# variable_delay_unit_1.tristate_inverter_1.en 0.11539f
C107 a_11340_352# en_4 6.99e-20
C108 en_1 en_0 0.010459f
C109 a_11340_772# variable_delay_unit_4.out 0.071074f
C110 en_3 variable_delay_unit_2.out 2.67e-19
C111 a_2496_352# a_2496_772# 0.011184f
C112 a_13406_352# variable_delay_unit_5.in 0.054206f
C113 variable_delay_unit_3.in variable_delay_unit_2.out 0.235667f
C114 variable_delay_unit_4.in a_14288_352# 7.65e-21
C115 a_7510_772# a_7510_352# 0.004142f
C116 variable_delay_unit_3.tristate_inverter_1.en a_10458_772# 0.11539f
C117 a_11340_772# a_11340_352# 0.011184f
C118 en_2 a_7510_772# 0.042718f
C119 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.out 0.085059f
C120 a_2496_772# in 7.65e-21
C121 a_8392_352# VDD 0.001468f
C122 VDD a_5444_772# 1.6584f
C123 a_1614_352# en_0 0.15982f
C124 a_4562_772# a_4562_352# 0.004142f
C125 variable_delay_unit_2.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en 0.002365f
C126 en_1 variable_delay_unit_2.out 0.043504f
C127 variable_delay_unit_3.tristate_inverter_1.en a_11340_352# 0.15982f
C128 variable_delay_unit_5.in en_4 0.574722f
C129 variable_delay_unit_3.out a_10458_352# 0.222585f
C130 VDD en_3 1.40792f
C131 variable_delay_unit_1.out a_5444_772# 0.493816f
C132 variable_delay_unit_3.in VDD 2.12807f
C133 a_2496_352# out 0.172055f
C134 VDD variable_delay_unit_4.in 2.12807f
C135 a_16354_352# VDD 0.160518f
C136 variable_delay_unit_3.out variable_delay_unit_2.out 0.071795f
C137 out in 0.487038f
C138 a_8392_772# variable_delay_unit_2.tristate_inverter_1.en 0.029284f
C139 variable_delay_unit_1.in VDD 2.12798f
C140 VDD en_1 1.40792f
C141 a_17236_772# variable_delay_unit_5.in 7.65e-21
C142 variable_delay_unit_5.in variable_delay_unit_3.tristate_inverter_1.en 7.91e-21
C143 variable_delay_unit_1.in variable_delay_unit_1.out 0.499092f
C144 a_2496_772# out 0.493816f
C145 a_14288_352# en_4 0.001909f
C146 a_13406_352# VDD 6.98e-19
C147 variable_delay_unit_1.out en_1 0.224474f
C148 VDD variable_delay_unit_3.out 1.34424f
C149 out variable_delay_unit_1.tristate_inverter_1.en 0.002141f
C150 VDD a_1614_352# 6.98e-19
C151 a_14288_772# variable_delay_unit_5.out 0.071074f
C152 a_4562_352# variable_delay_unit_1.tristate_inverter_1.en 2.39e-19
C153 a_10458_352# variable_delay_unit_3.tristate_inverter_1.en 2.39e-19
C154 a_8392_352# variable_delay_unit_2.in 7.65e-21
C155 variable_delay_unit_2.in a_5444_772# 0.020173f
C156 a_1614_772# variable_delay_unit_0.tristate_inverter_1.en 0.11539f
C157 VDD en_4 1.41838f
C158 variable_delay_unit_5.forward variable_delay_unit_5.tristate_inverter_1.en 0.794183f
C159 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_2.out 0.002141f
C160 variable_delay_unit_3.in variable_delay_unit_2.in 0.087283f
C161 VDD a_11340_772# 1.6584f
C162 variable_delay_unit_5.forward variable_delay_unit_5.out 0.234428f
C163 variable_delay_unit_1.in variable_delay_unit_2.in 0.087283f
C164 a_5444_352# a_5444_772# 0.011184f
C165 VDD a_17236_772# 1.78268f
C166 variable_delay_unit_2.in en_1 0.574722f
C167 VDD variable_delay_unit_3.tristate_inverter_1.en 2.77611f
C168 variable_delay_unit_1.in a_5444_352# 7.65e-21
C169 variable_delay_unit_1.in a_4562_772# 8.82e-20
C170 variable_delay_unit_4.out variable_delay_unit_4.tristate_inverter_1.en 0.12029f
C171 a_8392_352# variable_delay_unit_2.tristate_inverter_1.en 0.15982f
C172 a_5444_352# en_1 0.001909f
C173 en_1 a_4562_772# 0.042718f
C174 variable_delay_unit_5.tristate_inverter_1.en variable_delay_unit_5.out 0.12029f
C175 a_14288_772# variable_delay_unit_4.in 7.65e-21
C176 en_3 variable_delay_unit_2.tristate_inverter_1.en 9.38e-20
C177 variable_delay_unit_3.in variable_delay_unit_2.tristate_inverter_1.en 0.814958f
C178 variable_delay_unit_4.in variable_delay_unit_2.tristate_inverter_1.en 7.91e-21
C179 variable_delay_unit_2.out a_7510_352# 0.222585f
C180 en_2 variable_delay_unit_2.out 0.224474f
C181 a_2496_352# en_1 6.99e-20
C182 a_5444_772# variable_delay_unit_1.tristate_inverter_1.en 0.029284f
C183 variable_delay_unit_1.in in 0.08442f
C184 en_1 variable_delay_unit_2.tristate_inverter_1.en 1.5e-19
C185 variable_delay_unit_3.in variable_delay_unit_1.tristate_inverter_1.en 7.91e-21
C186 a_17236_352# variable_delay_unit_5.in 7.65e-21
C187 a_16354_352# variable_delay_unit_5.forward 0.054206f
C188 variable_delay_unit_5.in variable_delay_unit_4.tristate_inverter_1.en 0.814958f
C189 VDD a_7510_352# 6.98e-19
C190 variable_delay_unit_1.in a_2496_772# 0.020173f
C191 a_8392_352# a_8392_772# 0.011184f
C192 VDD en_2 1.40792f
C193 a_2496_772# en_1 6.99e-20
C194 en_0 variable_delay_unit_0.tristate_inverter_1.en 1.09349f
C195 variable_delay_unit_3.out variable_delay_unit_2.tristate_inverter_1.en 0.085059f
C196 variable_delay_unit_1.in variable_delay_unit_1.tristate_inverter_1.en 0.09141f
C197 en_3 a_8392_772# 6.99e-20
C198 variable_delay_unit_3.in a_8392_772# 0.020173f
C199 en_2 variable_delay_unit_1.out 2.67e-19
C200 en_1 variable_delay_unit_1.tristate_inverter_1.en 1.09349f
C201 a_1614_352# in 8.82e-20
C202 a_14288_772# en_4 0.124274f
C203 variable_delay_unit_1.in out 0.235655f
C204 a_1614_772# en_0 0.042718f
C205 variable_delay_unit_4.tristate_inverter_1.en a_14288_352# 0.15982f
C206 out en_1 2.67e-19
C207 variable_delay_unit_1.in a_4562_352# 8.82e-20
C208 a_16354_352# variable_delay_unit_5.tristate_inverter_1.en 2.39e-19
C209 variable_delay_unit_2.out a_7510_772# 0.505512f
C210 a_13406_772# variable_delay_unit_4.in 8.82e-20
C211 en_1 a_4562_352# 0.15982f
C212 variable_delay_unit_5.forward en_4 3.37e-20
C213 variable_delay_unit_3.out a_8392_772# 0.071074f
C214 a_11340_352# variable_delay_unit_4.out 0.070146f
C215 a_17236_352# VDD 0.003377f
C216 VDD variable_delay_unit_4.tristate_inverter_1.en 2.7762f
C217 a_16354_352# variable_delay_unit_5.out 0.222585f
C218 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_2.tristate_inverter_1.en 0.002365f
C219 variable_delay_unit_2.in a_7510_352# 8.82e-20
C220 out a_1614_352# 0.222585f
C221 VDD variable_delay_unit_0.tristate_inverter_1.en 2.77513f
C222 variable_delay_unit_2.in en_2 0.506369f
C223 VDD a_7510_772# 1.6584f
C224 a_17236_772# variable_delay_unit_5.forward 0.016896f
C225 variable_delay_unit_1.out variable_delay_unit_0.tristate_inverter_1.en 0.085059f
C226 a_13406_352# a_13406_772# 0.004142f
C227 variable_delay_unit_5.in variable_delay_unit_4.out 0.235667f
C228 VDD a_1614_772# 1.6584f
C229 a_16354_772# variable_delay_unit_5.in 8.82e-20
C230 a_5444_352# en_2 6.99e-20
C231 en_4 variable_delay_unit_5.tristate_inverter_1.en 1.5e-19
C232 a_10458_352# a_10458_772# 0.004142f
C233 a_13406_772# en_4 0.042718f
C234 en_4 variable_delay_unit_5.out 0.043504f
C235 a_8392_352# en_3 6.99e-20
C236 variable_delay_unit_4.out a_14288_352# 0.172055f
C237 a_17236_772# variable_delay_unit_5.tristate_inverter_1.en 0.029284f
C238 a_7510_352# variable_delay_unit_2.tristate_inverter_1.en 2.39e-19
C239 variable_delay_unit_3.in en_3 0.506369f
C240 variable_delay_unit_2.in variable_delay_unit_0.tristate_inverter_1.en 7.91e-21
C241 en_3 variable_delay_unit_4.in 0.574722f
C242 en_2 variable_delay_unit_2.tristate_inverter_1.en 1.09349f
C243 variable_delay_unit_1.in a_5444_772# 7.65e-21
C244 variable_delay_unit_3.in variable_delay_unit_4.in 0.087283f
C245 variable_delay_unit_2.in a_7510_772# 8.82e-20
C246 en_1 a_5444_772# 0.124274f
C247 a_17236_772# variable_delay_unit_5.out 0.493816f
C248 VDD a_10458_772# 1.6584f
C249 VDD variable_delay_unit_4.out 1.3445f
C250 variable_delay_unit_3.in en_1 3.37e-20
C251 a_8392_352# variable_delay_unit_3.out 0.070146f
C252 VDD a_16354_772# 1.70112f
C253 en_2 variable_delay_unit_1.tristate_inverter_1.en 9.38e-20
C254 VDD a_11340_352# 0.001468f
C255 variable_delay_unit_1.in en_1 0.506369f
C256 en_3 variable_delay_unit_3.out 0.224474f
C257 a_13406_352# variable_delay_unit_4.in 8.82e-20
C258 variable_delay_unit_3.in variable_delay_unit_3.out 0.499092f
C259 variable_delay_unit_3.out variable_delay_unit_4.in 0.235667f
C260 en_2 a_8392_772# 0.124274f
C261 a_2496_352# variable_delay_unit_0.tristate_inverter_1.en 0.15982f
C262 a_14288_772# variable_delay_unit_4.tristate_inverter_1.en 0.029284f
C263 en_3 en_4 0.010459f
C264 variable_delay_unit_4.in en_4 0.506369f
C265 VDD variable_delay_unit_5.in 2.63444f
C266 variable_delay_unit_1.in a_1614_352# 0.054206f
C267 in variable_delay_unit_0.tristate_inverter_1.en 0.091118f
C268 VDD en_0 1.41013f
C269 a_11340_772# en_3 0.124274f
C270 a_7510_772# variable_delay_unit_2.tristate_inverter_1.en 0.11539f
C271 variable_delay_unit_3.in a_11340_772# 7.65e-21
C272 a_11340_772# variable_delay_unit_4.in 0.020173f
C273 a_2496_772# variable_delay_unit_0.tristate_inverter_1.en 0.029284f
C274 variable_delay_unit_5.forward variable_delay_unit_4.tristate_inverter_1.en 7.91e-21
C275 variable_delay_unit_1.out en_0 0.043504f
C276 VDD a_10458_352# 6.98e-19
C277 a_1614_772# in 8.82e-20
C278 en_3 variable_delay_unit_3.tristate_inverter_1.en 1.09349f
C279 variable_delay_unit_0.tristate_inverter_1.en variable_delay_unit_1.tristate_inverter_1.en 0.002365f
C280 variable_delay_unit_3.in variable_delay_unit_3.tristate_inverter_1.en 0.09141f
C281 variable_delay_unit_3.tristate_inverter_1.en variable_delay_unit_4.in 0.814958f
C282 a_13406_352# en_4 0.15982f
C283 variable_delay_unit_3.out en_4 2.67e-19
C284 VDD variable_delay_unit_2.out 1.34424f
C285 VDD a_14288_352# 0.001538f
C286 out variable_delay_unit_0.tristate_inverter_1.en 0.12022f
C287 a_11340_772# variable_delay_unit_3.out 0.493816f
C288 variable_delay_unit_1.out variable_delay_unit_2.out 0.071795f
C289 variable_delay_unit_3.out variable_delay_unit_3.tristate_inverter_1.en 0.12029f
C290 a_17236_352# variable_delay_unit_5.tristate_inverter_1.en 0.15982f
C291 variable_delay_unit_4.tristate_inverter_1.en variable_delay_unit_5.tristate_inverter_1.en 0.002365f
C292 a_11340_772# en_4 6.99e-20
C293 variable_delay_unit_2.in en_0 3.37e-20
C294 out a_1614_772# 0.505512f
C295 a_13406_772# variable_delay_unit_4.tristate_inverter_1.en 0.11539f
C296 en_4 VSS 2.08969f
C297 en_3 VSS 2.08969f
C298 en_2 VSS 2.08969f
C299 en_1 VSS 2.08969f
C300 out VSS 1.89289f
C301 in VSS 1.0591f
C302 en_0 VSS 2.22578f
C303 VDD VSS 52.60628f
C304 a_17236_352# VSS 0.784074f
C305 a_16354_352# VSS 0.71648f
C306 a_14288_352# VSS 0.717347f
C307 a_13406_352# VSS 0.71648f
C308 a_17236_772# VSS 0.114203f
C309 a_16354_772# VSS 0.037888f
C310 variable_delay_unit_5.forward VSS 2.632682f
C311 variable_delay_unit_5.tristate_inverter_1.en VSS 2.962361f
C312 a_11340_352# VSS 0.717347f
C313 a_10458_352# VSS 0.71648f
C314 a_14288_772# VSS 0.043128f
C315 variable_delay_unit_5.out VSS 2.29732f
C316 a_13406_772# VSS 0.037888f
C317 variable_delay_unit_5.in VSS 3.857309f
C318 variable_delay_unit_4.tristate_inverter_1.en VSS 2.51692f
C319 a_8392_352# VSS 0.717347f
C320 a_7510_352# VSS 0.71648f
C321 a_11340_772# VSS 0.043128f
C322 variable_delay_unit_4.out VSS 2.21957f
C323 a_10458_772# VSS 0.037888f
C324 variable_delay_unit_4.in VSS 3.60152f
C325 variable_delay_unit_3.tristate_inverter_1.en VSS 2.51692f
C326 a_5444_352# VSS 0.717347f
C327 a_4562_352# VSS 0.71648f
C328 a_8392_772# VSS 0.043128f
C329 variable_delay_unit_3.out VSS 2.21957f
C330 a_7510_772# VSS 0.037888f
C331 variable_delay_unit_3.in VSS 3.60152f
C332 variable_delay_unit_2.tristate_inverter_1.en VSS 2.51692f
C333 a_2496_352# VSS 0.717347f
C334 a_1614_352# VSS 0.71648f
C335 a_5444_772# VSS 0.043128f
C336 variable_delay_unit_2.out VSS 2.21957f
C337 a_4562_772# VSS 0.037888f
C338 variable_delay_unit_2.in VSS 3.60152f
C339 variable_delay_unit_1.tristate_inverter_1.en VSS 2.51692f
C340 a_2496_772# VSS 0.043128f
C341 variable_delay_unit_1.out VSS 2.21957f
C342 a_1614_772# VSS 0.037888f
C343 variable_delay_unit_1.in VSS 3.60479f
C344 variable_delay_unit_0.tristate_inverter_1.en VSS 2.52279f
C345 variable_delay_unit_3.tristate_inverter_1.en.t4 VSS 0.019446f
C346 variable_delay_unit_3.tristate_inverter_1.en.t2 VSS 0.025128f
C347 variable_delay_unit_3.tristate_inverter_1.en.t7 VSS 0.025128f
C348 variable_delay_unit_3.tristate_inverter_1.en.n0 VSS 0.074066f
C349 variable_delay_unit_3.tristate_inverter_1.en.t1 VSS 0.154367f
C350 variable_delay_unit_3.tristate_inverter_1.en.t0 VSS 0.048564f
C351 variable_delay_unit_3.tristate_inverter_1.en.n1 VSS 0.616703f
C352 variable_delay_unit_3.tristate_inverter_1.en.n2 VSS 0.678061f
C353 variable_delay_unit_3.tristate_inverter_1.en.t6 VSS 0.066961f
C354 variable_delay_unit_3.tristate_inverter_1.en.t3 VSS 0.062029f
C355 variable_delay_unit_3.tristate_inverter_1.en.t5 VSS 0.067187f
C356 variable_delay_unit_3.tristate_inverter_1.en.n3 VSS 0.065756f
C357 variable_delay_unit_3.tristate_inverter_1.en.n4 VSS 0.045654f
C358 variable_delay_unit_4.tristate_inverter_1.en.t6 VSS 0.019446f
C359 variable_delay_unit_4.tristate_inverter_1.en.t4 VSS 0.025128f
C360 variable_delay_unit_4.tristate_inverter_1.en.t2 VSS 0.025128f
C361 variable_delay_unit_4.tristate_inverter_1.en.n0 VSS 0.074066f
C362 variable_delay_unit_4.tristate_inverter_1.en.t1 VSS 0.154367f
C363 variable_delay_unit_4.tristate_inverter_1.en.t0 VSS 0.048564f
C364 variable_delay_unit_4.tristate_inverter_1.en.n1 VSS 0.616703f
C365 variable_delay_unit_4.tristate_inverter_1.en.n2 VSS 0.678061f
C366 variable_delay_unit_4.tristate_inverter_1.en.t7 VSS 0.066961f
C367 variable_delay_unit_4.tristate_inverter_1.en.t3 VSS 0.062029f
C368 variable_delay_unit_4.tristate_inverter_1.en.t5 VSS 0.067187f
C369 variable_delay_unit_4.tristate_inverter_1.en.n3 VSS 0.065756f
C370 variable_delay_unit_4.tristate_inverter_1.en.n4 VSS 0.045654f
C371 variable_delay_unit_1.in.t2 VSS 0.044984f
C372 variable_delay_unit_1.in.t3 VSS 0.017058f
C373 variable_delay_unit_1.in.n0 VSS 0.04731f
C374 variable_delay_unit_1.in.t1 VSS 0.033139f
C375 variable_delay_unit_1.in.t0 VSS 0.105354f
C376 variable_delay_unit_1.in.n1 VSS 0.255341f
C377 variable_delay_unit_1.in.t4 VSS 0.042943f
C378 variable_delay_unit_1.in.t5 VSS 0.013862f
C379 variable_delay_unit_1.in.n2 VSS 0.045159f
C380 variable_delay_unit_1.in.n3 VSS 0.420531f
C381 variable_delay_unit_5.forward.t2 VSS 0.067654f
C382 variable_delay_unit_5.forward.t3 VSS 0.025654f
C383 variable_delay_unit_5.forward.n0 VSS 0.071153f
C384 variable_delay_unit_5.forward.t0 VSS 0.04984f
C385 variable_delay_unit_5.forward.t1 VSS 0.15845f
C386 variable_delay_unit_5.forward.n1 VSS 0.384027f
C387 variable_delay_unit_5.forward.n2 VSS 0.632469f
C388 variable_delay_unit_5.in.t4 VSS 0.055694f
C389 variable_delay_unit_5.in.t5 VSS 0.021119f
C390 variable_delay_unit_5.in.n0 VSS 0.058574f
C391 variable_delay_unit_5.in.t0 VSS 0.041029f
C392 variable_delay_unit_5.in.t1 VSS 0.130438f
C393 variable_delay_unit_5.in.n1 VSS 0.316137f
C394 variable_delay_unit_5.in.t2 VSS 0.053167f
C395 variable_delay_unit_5.in.t3 VSS 0.017162f
C396 variable_delay_unit_5.in.n2 VSS 0.055911f
C397 variable_delay_unit_5.in.n3 VSS 0.520657f
C398 variable_delay_unit_0.tristate_inverter_1.en.t4 VSS 0.019446f
C399 variable_delay_unit_0.tristate_inverter_1.en.t2 VSS 0.025128f
C400 variable_delay_unit_0.tristate_inverter_1.en.t6 VSS 0.025128f
C401 variable_delay_unit_0.tristate_inverter_1.en.n0 VSS 0.074066f
C402 variable_delay_unit_0.tristate_inverter_1.en.t1 VSS 0.154367f
C403 variable_delay_unit_0.tristate_inverter_1.en.t0 VSS 0.048564f
C404 variable_delay_unit_0.tristate_inverter_1.en.n1 VSS 0.616703f
C405 variable_delay_unit_0.tristate_inverter_1.en.n2 VSS 0.678061f
C406 variable_delay_unit_0.tristate_inverter_1.en.t5 VSS 0.066961f
C407 variable_delay_unit_0.tristate_inverter_1.en.t7 VSS 0.062029f
C408 variable_delay_unit_0.tristate_inverter_1.en.t3 VSS 0.067187f
C409 variable_delay_unit_0.tristate_inverter_1.en.n3 VSS 0.065756f
C410 variable_delay_unit_0.tristate_inverter_1.en.n4 VSS 0.045654f
C411 variable_delay_unit_1.tristate_inverter_1.en.t5 VSS 0.019446f
C412 variable_delay_unit_1.tristate_inverter_1.en.t2 VSS 0.025128f
C413 variable_delay_unit_1.tristate_inverter_1.en.t3 VSS 0.025128f
C414 variable_delay_unit_1.tristate_inverter_1.en.n0 VSS 0.074066f
C415 variable_delay_unit_1.tristate_inverter_1.en.t1 VSS 0.154367f
C416 variable_delay_unit_1.tristate_inverter_1.en.t0 VSS 0.048564f
C417 variable_delay_unit_1.tristate_inverter_1.en.n1 VSS 0.616703f
C418 variable_delay_unit_1.tristate_inverter_1.en.n2 VSS 0.678061f
C419 variable_delay_unit_1.tristate_inverter_1.en.t7 VSS 0.066961f
C420 variable_delay_unit_1.tristate_inverter_1.en.t4 VSS 0.062029f
C421 variable_delay_unit_1.tristate_inverter_1.en.t6 VSS 0.067187f
C422 variable_delay_unit_1.tristate_inverter_1.en.n3 VSS 0.065756f
C423 variable_delay_unit_1.tristate_inverter_1.en.n4 VSS 0.045654f
C424 variable_delay_unit_2.in.t4 VSS 0.044984f
C425 variable_delay_unit_2.in.t5 VSS 0.017058f
C426 variable_delay_unit_2.in.n0 VSS 0.04731f
C427 variable_delay_unit_2.in.t1 VSS 0.033139f
C428 variable_delay_unit_2.in.t0 VSS 0.105354f
C429 variable_delay_unit_2.in.n1 VSS 0.255341f
C430 variable_delay_unit_2.in.t2 VSS 0.042943f
C431 variable_delay_unit_2.in.t3 VSS 0.013862f
C432 variable_delay_unit_2.in.n2 VSS 0.045159f
C433 variable_delay_unit_2.in.n3 VSS 0.420531f
C434 variable_delay_unit_4.in.t3 VSS 0.044984f
C435 variable_delay_unit_4.in.t5 VSS 0.017058f
C436 variable_delay_unit_4.in.n0 VSS 0.04731f
C437 variable_delay_unit_4.in.t0 VSS 0.033139f
C438 variable_delay_unit_4.in.t1 VSS 0.105354f
C439 variable_delay_unit_4.in.n1 VSS 0.255341f
C440 variable_delay_unit_4.in.t2 VSS 0.042943f
C441 variable_delay_unit_4.in.t4 VSS 0.013862f
C442 variable_delay_unit_4.in.n2 VSS 0.045159f
C443 variable_delay_unit_4.in.n3 VSS 0.420531f
C444 variable_delay_unit_3.in.t4 VSS 0.044984f
C445 variable_delay_unit_3.in.t5 VSS 0.017058f
C446 variable_delay_unit_3.in.n0 VSS 0.04731f
C447 variable_delay_unit_3.in.t0 VSS 0.033139f
C448 variable_delay_unit_3.in.t1 VSS 0.105354f
C449 variable_delay_unit_3.in.n1 VSS 0.255341f
C450 variable_delay_unit_3.in.t2 VSS 0.042943f
C451 variable_delay_unit_3.in.t3 VSS 0.013862f
C452 variable_delay_unit_3.in.n2 VSS 0.045159f
C453 variable_delay_unit_3.in.n3 VSS 0.420531f
C454 variable_delay_unit_2.tristate_inverter_1.en.t6 VSS 0.019446f
C455 variable_delay_unit_2.tristate_inverter_1.en.t4 VSS 0.025128f
C456 variable_delay_unit_2.tristate_inverter_1.en.t2 VSS 0.025128f
C457 variable_delay_unit_2.tristate_inverter_1.en.n0 VSS 0.074066f
C458 variable_delay_unit_2.tristate_inverter_1.en.t0 VSS 0.154367f
C459 variable_delay_unit_2.tristate_inverter_1.en.t1 VSS 0.048564f
C460 variable_delay_unit_2.tristate_inverter_1.en.n1 VSS 0.616703f
C461 variable_delay_unit_2.tristate_inverter_1.en.n2 VSS 0.678061f
C462 variable_delay_unit_2.tristate_inverter_1.en.t7 VSS 0.066961f
C463 variable_delay_unit_2.tristate_inverter_1.en.t3 VSS 0.062029f
C464 variable_delay_unit_2.tristate_inverter_1.en.t5 VSS 0.067187f
C465 variable_delay_unit_2.tristate_inverter_1.en.n3 VSS 0.065756f
C466 variable_delay_unit_2.tristate_inverter_1.en.n4 VSS 0.045654f
C467 VDD.n0 VSS 0.167082f
C468 VDD.t12 VSS 0.04115f
C469 VDD.n1 VSS 0.042641f
C470 VDD.n2 VSS 0.038087f
C471 VDD.n3 VSS 0.025131f
C472 VDD.t101 VSS 0.171896f
C473 VDD.n4 VSS 0.049621f
C474 VDD.n5 VSS 0.049621f
C475 VDD.t102 VSS 0.04115f
C476 VDD.n6 VSS 0.017155f
C477 VDD.n7 VSS 0.167082f
C478 VDD.n8 VSS 0.046707f
C479 VDD.t22 VSS 0.010965f
C480 VDD.t108 VSS 0.010965f
C481 VDD.n9 VSS 0.032003f
C482 VDD.t46 VSS 0.040485f
C483 VDD.n10 VSS 0.14597f
C484 VDD.n11 VSS 0.063111f
C485 VDD.n12 VSS 0.046707f
C486 VDD.n13 VSS 0.029558f
C487 VDD.n14 VSS 0.161197f
C488 VDD.t106 VSS 0.137724f
C489 VDD.n15 VSS 0.076238f
C490 VDD.n16 VSS 0.076238f
C491 VDD.t14 VSS 0.010965f
C492 VDD.t24 VSS 0.010965f
C493 VDD.n17 VSS 0.032003f
C494 VDD.t54 VSS 0.040485f
C495 VDD.n18 VSS 0.14597f
C496 VDD.t23 VSS 0.07836f
C497 VDD.n19 VSS 0.05224f
C498 VDD.t13 VSS 0.07836f
C499 VDD.t53 VSS 0.154493f
C500 VDD.n20 VSS 0.161197f
C501 VDD.n21 VSS 0.046707f
C502 VDD.n22 VSS 0.167082f
C503 VDD.t33 VSS 0.04115f
C504 VDD.n23 VSS 0.042641f
C505 VDD.n24 VSS 0.038087f
C506 VDD.n25 VSS 0.025131f
C507 VDD.t39 VSS 0.171896f
C508 VDD.n26 VSS 0.049621f
C509 VDD.n27 VSS 0.049621f
C510 VDD.t40 VSS 0.04115f
C511 VDD.n28 VSS 0.017155f
C512 VDD.n29 VSS 0.167082f
C513 VDD.n30 VSS 0.046707f
C514 VDD.t38 VSS 0.010965f
C515 VDD.t94 VSS 0.010965f
C516 VDD.n31 VSS 0.032003f
C517 VDD.t92 VSS 0.040485f
C518 VDD.n32 VSS 0.14597f
C519 VDD.n33 VSS 0.063111f
C520 VDD.n34 VSS 0.046707f
C521 VDD.n35 VSS 0.029558f
C522 VDD.n36 VSS 0.161197f
C523 VDD.t104 VSS 0.137724f
C524 VDD.n37 VSS 0.076238f
C525 VDD.n38 VSS 0.076238f
C526 VDD.t42 VSS 0.010965f
C527 VDD.t88 VSS 0.010965f
C528 VDD.n39 VSS 0.032003f
C529 VDD.t20 VSS 0.040485f
C530 VDD.n40 VSS 0.14597f
C531 VDD.t87 VSS 0.07836f
C532 VDD.n41 VSS 0.05224f
C533 VDD.t41 VSS 0.07836f
C534 VDD.t19 VSS 0.154493f
C535 VDD.n42 VSS 0.161197f
C536 VDD.n43 VSS 0.046707f
C537 VDD.n44 VSS 0.167082f
C538 VDD.t59 VSS 0.04115f
C539 VDD.n45 VSS 0.042641f
C540 VDD.n46 VSS 0.038087f
C541 VDD.n47 VSS 0.025131f
C542 VDD.t3 VSS 0.171896f
C543 VDD.n48 VSS 0.049621f
C544 VDD.n49 VSS 0.049621f
C545 VDD.t4 VSS 0.04115f
C546 VDD.n50 VSS 0.017155f
C547 VDD.n51 VSS 0.167082f
C548 VDD.n52 VSS 0.046707f
C549 VDD.t64 VSS 0.010965f
C550 VDD.t66 VSS 0.010965f
C551 VDD.n53 VSS 0.032003f
C552 VDD.t98 VSS 0.040485f
C553 VDD.n54 VSS 0.14597f
C554 VDD.n55 VSS 0.063111f
C555 VDD.n56 VSS 0.046707f
C556 VDD.n57 VSS 0.029558f
C557 VDD.n58 VSS 0.161197f
C558 VDD.t105 VSS 0.137724f
C559 VDD.n59 VSS 0.076238f
C560 VDD.n60 VSS 0.076238f
C561 VDD.t10 VSS 0.010965f
C562 VDD.t16 VSS 0.010965f
C563 VDD.n61 VSS 0.032003f
C564 VDD.t52 VSS 0.040485f
C565 VDD.n62 VSS 0.14597f
C566 VDD.t15 VSS 0.07836f
C567 VDD.n63 VSS 0.05224f
C568 VDD.t9 VSS 0.07836f
C569 VDD.t51 VSS 0.154493f
C570 VDD.n64 VSS 0.161197f
C571 VDD.n65 VSS 0.046707f
C572 VDD.n66 VSS 0.167082f
C573 VDD.t2 VSS 0.04115f
C574 VDD.n67 VSS 0.042641f
C575 VDD.n68 VSS 0.038087f
C576 VDD.n69 VSS 0.025131f
C577 VDD.t109 VSS 0.171896f
C578 VDD.n70 VSS 0.049621f
C579 VDD.n71 VSS 0.049621f
C580 VDD.t110 VSS 0.04115f
C581 VDD.n72 VSS 0.017155f
C582 VDD.n73 VSS 0.167082f
C583 VDD.n74 VSS 0.046707f
C584 VDD.t62 VSS 0.010965f
C585 VDD.t18 VSS 0.010965f
C586 VDD.n75 VSS 0.032003f
C587 VDD.t8 VSS 0.040485f
C588 VDD.n76 VSS 0.14597f
C589 VDD.n77 VSS 0.063111f
C590 VDD.n78 VSS 0.046707f
C591 VDD.n79 VSS 0.029558f
C592 VDD.n80 VSS 0.161197f
C593 VDD.t103 VSS 0.137724f
C594 VDD.n81 VSS 0.076238f
C595 VDD.n82 VSS 0.076238f
C596 VDD.t44 VSS 0.010965f
C597 VDD.t57 VSS 0.010965f
C598 VDD.n83 VSS 0.032003f
C599 VDD.t30 VSS 0.040485f
C600 VDD.n84 VSS 0.14597f
C601 VDD.t56 VSS 0.07836f
C602 VDD.n85 VSS 0.05224f
C603 VDD.t43 VSS 0.07836f
C604 VDD.t29 VSS 0.154493f
C605 VDD.n86 VSS 0.161197f
C606 VDD.n87 VSS 0.046707f
C607 VDD.n88 VSS 0.167082f
C608 VDD.t71 VSS 0.04115f
C609 VDD.n89 VSS 0.042641f
C610 VDD.n90 VSS 0.038087f
C611 VDD.n91 VSS 0.025131f
C612 VDD.t95 VSS 0.171896f
C613 VDD.n92 VSS 0.049621f
C614 VDD.n93 VSS 0.049621f
C615 VDD.t96 VSS 0.04115f
C616 VDD.n94 VSS 0.017155f
C617 VDD.n95 VSS 0.167082f
C618 VDD.n96 VSS 0.046707f
C619 VDD.t86 VSS 0.010965f
C620 VDD.t84 VSS 0.010965f
C621 VDD.n97 VSS 0.032003f
C622 VDD.t82 VSS 0.040485f
C623 VDD.n98 VSS 0.14597f
C624 VDD.n99 VSS 0.063111f
C625 VDD.n100 VSS 0.046707f
C626 VDD.n101 VSS 0.029558f
C627 VDD.n102 VSS 0.161197f
C628 VDD.t36 VSS 0.137724f
C629 VDD.n103 VSS 0.076238f
C630 VDD.n104 VSS 0.076238f
C631 VDD.t74 VSS 0.010965f
C632 VDD.t80 VSS 0.010965f
C633 VDD.n105 VSS 0.032003f
C634 VDD.t77 VSS 0.040485f
C635 VDD.n106 VSS 0.14597f
C636 VDD.t79 VSS 0.07836f
C637 VDD.n107 VSS 0.05224f
C638 VDD.t73 VSS 0.07836f
C639 VDD.t76 VSS 0.154493f
C640 VDD.n108 VSS 0.161197f
C641 VDD.n109 VSS 0.046817f
C642 VDD.n110 VSS 0.029382f
C643 VDD.n111 VSS 0.027345f
C644 VDD.n112 VSS 0.063111f
C645 VDD.n113 VSS 0.046707f
C646 VDD.n114 VSS 0.029558f
C647 VDD.n115 VSS 0.281383f
C648 VDD.n116 VSS 0.281383f
C649 VDD.t31 VSS 0.137724f
C650 VDD.t85 VSS 0.07836f
C651 VDD.t81 VSS 0.154493f
C652 VDD.t83 VSS 0.07836f
C653 VDD.n117 VSS 0.05224f
C654 VDD.n118 VSS 0.076238f
C655 VDD.n119 VSS 0.076238f
C656 VDD.n120 VSS 0.027345f
C657 VDD.n121 VSS 0.029684f
C658 VDD.n122 VSS 0.035706f
C659 VDD.n123 VSS 0.059342f
C660 VDD.n124 VSS 0.011434f
C661 VDD.n125 VSS 0.075919f
C662 VDD.n126 VSS 0.039979f
C663 VDD.n127 VSS 0.038087f
C664 VDD.n128 VSS 0.025131f
C665 VDD.n129 VSS 0.136478f
C666 VDD.n130 VSS 0.136478f
C667 VDD.t70 VSS 0.171896f
C668 VDD.n131 VSS 0.017155f
C669 VDD.n132 VSS 0.049621f
C670 VDD.n133 VSS 0.049621f
C671 VDD.n134 VSS 0.011434f
C672 VDD.n135 VSS 0.075919f
C673 VDD.n136 VSS 0.041776f
C674 VDD.t113 VSS 0.00518f
C675 VDD.t112 VSS 0.006694f
C676 VDD.t115 VSS 0.006694f
C677 VDD.n137 VSS 0.01973f
C678 VDD.t72 VSS 0.016524f
C679 VDD.t75 VSS 0.017898f
C680 VDD.n138 VSS 0.017516f
C681 VDD.t78 VSS 0.017838f
C682 VDD.n139 VSS 0.012162f
C683 VDD.n140 VSS 0.127782f
C684 VDD.n141 VSS 0.100401f
C685 VDD.t69 VSS 0.01675f
C686 VDD.t114 VSS 0.005407f
C687 VDD.n142 VSS 0.01651f
C688 VDD.n143 VSS 0.118699f
C689 VDD.n144 VSS 0.037504f
C690 VDD.n145 VSS 0.029958f
C691 VDD.n146 VSS 0.029382f
C692 VDD.n147 VSS 0.027345f
C693 VDD.n148 VSS 0.063111f
C694 VDD.n149 VSS 0.046707f
C695 VDD.n150 VSS 0.029558f
C696 VDD.n151 VSS 0.281383f
C697 VDD.n152 VSS 0.281383f
C698 VDD.t55 VSS 0.137724f
C699 VDD.t61 VSS 0.07836f
C700 VDD.t7 VSS 0.154493f
C701 VDD.t17 VSS 0.07836f
C702 VDD.n153 VSS 0.05224f
C703 VDD.n154 VSS 0.076238f
C704 VDD.n155 VSS 0.076238f
C705 VDD.n156 VSS 0.027345f
C706 VDD.n157 VSS 0.029684f
C707 VDD.n158 VSS 0.035706f
C708 VDD.n159 VSS 0.059342f
C709 VDD.n160 VSS 0.011434f
C710 VDD.n161 VSS 0.075919f
C711 VDD.n162 VSS 0.039979f
C712 VDD.n163 VSS 0.038087f
C713 VDD.n164 VSS 0.025131f
C714 VDD.n165 VSS 0.136478f
C715 VDD.n166 VSS 0.136478f
C716 VDD.t1 VSS 0.171896f
C717 VDD.n167 VSS 0.017155f
C718 VDD.n168 VSS 0.049621f
C719 VDD.n169 VSS 0.049621f
C720 VDD.n170 VSS 0.011434f
C721 VDD.n171 VSS 0.075919f
C722 VDD.n172 VSS 0.067496f
C723 VDD.n173 VSS 0.029958f
C724 VDD.n174 VSS 0.029382f
C725 VDD.n175 VSS 0.027345f
C726 VDD.n176 VSS 0.063111f
C727 VDD.n177 VSS 0.046707f
C728 VDD.n178 VSS 0.029558f
C729 VDD.n179 VSS 0.281383f
C730 VDD.n180 VSS 0.281383f
C731 VDD.t111 VSS 0.137724f
C732 VDD.t63 VSS 0.07836f
C733 VDD.t97 VSS 0.154493f
C734 VDD.t65 VSS 0.07836f
C735 VDD.n181 VSS 0.05224f
C736 VDD.n182 VSS 0.076238f
C737 VDD.n183 VSS 0.076238f
C738 VDD.n184 VSS 0.027345f
C739 VDD.n185 VSS 0.029684f
C740 VDD.n186 VSS 0.035706f
C741 VDD.n187 VSS 0.059342f
C742 VDD.n188 VSS 0.011434f
C743 VDD.n189 VSS 0.075919f
C744 VDD.n190 VSS 0.039979f
C745 VDD.n191 VSS 0.038087f
C746 VDD.n192 VSS 0.025131f
C747 VDD.n193 VSS 0.136478f
C748 VDD.n194 VSS 0.136478f
C749 VDD.t58 VSS 0.171896f
C750 VDD.n195 VSS 0.017155f
C751 VDD.n196 VSS 0.049621f
C752 VDD.n197 VSS 0.049621f
C753 VDD.n198 VSS 0.011434f
C754 VDD.n199 VSS 0.075919f
C755 VDD.n200 VSS 0.067496f
C756 VDD.n201 VSS 0.029958f
C757 VDD.n202 VSS 0.029382f
C758 VDD.n203 VSS 0.027345f
C759 VDD.n204 VSS 0.063111f
C760 VDD.n205 VSS 0.046707f
C761 VDD.n206 VSS 0.029558f
C762 VDD.n207 VSS 0.281383f
C763 VDD.n208 VSS 0.281383f
C764 VDD.t0 VSS 0.137724f
C765 VDD.t37 VSS 0.07836f
C766 VDD.t91 VSS 0.154493f
C767 VDD.t93 VSS 0.07836f
C768 VDD.n209 VSS 0.05224f
C769 VDD.n210 VSS 0.076238f
C770 VDD.n211 VSS 0.076238f
C771 VDD.n212 VSS 0.027345f
C772 VDD.n213 VSS 0.029684f
C773 VDD.n214 VSS 0.035706f
C774 VDD.n215 VSS 0.059342f
C775 VDD.n216 VSS 0.011434f
C776 VDD.n217 VSS 0.075919f
C777 VDD.n218 VSS 0.039979f
C778 VDD.n219 VSS 0.038087f
C779 VDD.n220 VSS 0.025131f
C780 VDD.n221 VSS 0.136478f
C781 VDD.n222 VSS 0.136478f
C782 VDD.t32 VSS 0.171896f
C783 VDD.n223 VSS 0.017155f
C784 VDD.n224 VSS 0.049621f
C785 VDD.n225 VSS 0.049621f
C786 VDD.n226 VSS 0.011434f
C787 VDD.n227 VSS 0.075919f
C788 VDD.n228 VSS 0.067496f
C789 VDD.n229 VSS 0.029958f
C790 VDD.n230 VSS 0.029382f
C791 VDD.n231 VSS 0.027345f
C792 VDD.n232 VSS 0.063111f
C793 VDD.n233 VSS 0.046707f
C794 VDD.n234 VSS 0.029558f
C795 VDD.n235 VSS 0.281383f
C796 VDD.n236 VSS 0.281383f
C797 VDD.t68 VSS 0.137724f
C798 VDD.t21 VSS 0.07836f
C799 VDD.t45 VSS 0.154493f
C800 VDD.t107 VSS 0.07836f
C801 VDD.n237 VSS 0.05224f
C802 VDD.n238 VSS 0.076238f
C803 VDD.n239 VSS 0.076238f
C804 VDD.n240 VSS 0.027345f
C805 VDD.n241 VSS 0.029684f
C806 VDD.n242 VSS 0.035706f
C807 VDD.n243 VSS 0.059342f
C808 VDD.n244 VSS 0.011434f
C809 VDD.n245 VSS 0.075919f
C810 VDD.n246 VSS 0.039979f
C811 VDD.n247 VSS 0.038087f
C812 VDD.n248 VSS 0.025131f
C813 VDD.n249 VSS 0.136478f
C814 VDD.n250 VSS 0.136478f
C815 VDD.t11 VSS 0.171896f
C816 VDD.n251 VSS 0.017155f
C817 VDD.n252 VSS 0.049621f
C818 VDD.n253 VSS 0.049621f
C819 VDD.n254 VSS 0.011434f
C820 VDD.n255 VSS 0.075919f
C821 VDD.n256 VSS 0.067496f
C822 VDD.n257 VSS 0.046707f
C823 VDD.t28 VSS 0.010965f
C824 VDD.t35 VSS 0.010965f
C825 VDD.n258 VSS 0.032003f
C826 VDD.t50 VSS 0.040485f
C827 VDD.n259 VSS 0.14597f
C828 VDD.n260 VSS 0.063111f
C829 VDD.n261 VSS 0.076238f
C830 VDD.n262 VSS 0.161197f
C831 VDD.t49 VSS 0.154493f
C832 VDD.t27 VSS 0.07836f
C833 VDD.n263 VSS 0.05224f
C834 VDD.t34 VSS 0.07836f
C835 VDD.t67 VSS 0.137724f
C836 VDD.t60 VSS 0.137724f
C837 VDD.n264 VSS 0.076238f
C838 VDD.n265 VSS 0.076238f
C839 VDD.t100 VSS 0.010965f
C840 VDD.t48 VSS 0.010965f
C841 VDD.n266 VSS 0.032003f
C842 VDD.t6 VSS 0.040485f
C843 VDD.n267 VSS 0.14597f
C844 VDD.t99 VSS 0.07836f
C845 VDD.n268 VSS 0.05224f
C846 VDD.t47 VSS 0.07836f
C847 VDD.t5 VSS 0.154493f
C848 VDD.n269 VSS 0.161197f
C849 VDD.n270 VSS 0.046707f
C850 VDD.n271 VSS 0.167082f
C851 VDD.t90 VSS 0.04115f
C852 VDD.n272 VSS 0.075919f
C853 VDD.n273 VSS 0.049621f
C854 VDD.n274 VSS 0.025131f
C855 VDD.n275 VSS 0.038087f
C856 VDD.t26 VSS 0.04115f
C857 VDD.n276 VSS 0.075919f
C858 VDD.n277 VSS 0.049621f
C859 VDD.n278 VSS 0.063382f
C860 VDD.n279 VSS 0.017155f
C861 VDD.t89 VSS 0.171896f
C862 VDD.n280 VSS 0.136478f
C863 VDD.n281 VSS 0.025131f
C864 VDD.n282 VSS 0.136478f
C865 VDD.t25 VSS 0.171896f
C866 VDD.n283 VSS 0.017155f
C867 VDD.n284 VSS 0.167082f
C868 VDD.n285 VSS 0.049621f
C869 VDD.n286 VSS 0.011434f
C870 VDD.n287 VSS 0.042641f
C871 VDD.n288 VSS 0.039979f
C872 VDD.n289 VSS 0.038087f
C873 VDD.n290 VSS 0.049621f
C874 VDD.n291 VSS 0.011434f
C875 VDD.n292 VSS 0.059342f
C876 VDD.n293 VSS 0.035706f
C877 VDD.n294 VSS 0.029684f
C878 VDD.n295 VSS 0.027345f
C879 VDD.n296 VSS 0.063111f
C880 VDD.n297 VSS 0.046707f
C881 VDD.n298 VSS 0.029558f
C882 VDD.n299 VSS 0.281383f
C883 VDD.n300 VSS 0.281383f
C884 VDD.n301 VSS 0.029558f
C885 VDD.n302 VSS 0.046707f
C886 VDD.n303 VSS 0.076238f
C887 VDD.n304 VSS 0.027345f
C888 VDD.n305 VSS 0.029382f
C889 VDD.n306 VSS 0.029958f
C890 variable_delay_unit_5.tristate_inverter_1.en.t6 VSS 0.027086f
C891 variable_delay_unit_5.tristate_inverter_1.en.t4 VSS 0.035f
C892 variable_delay_unit_5.tristate_inverter_1.en.t3 VSS 0.035f
C893 variable_delay_unit_5.tristate_inverter_1.en.n0 VSS 0.103163f
C894 variable_delay_unit_5.tristate_inverter_1.en.t1 VSS 0.215011f
C895 variable_delay_unit_5.tristate_inverter_1.en.t0 VSS 0.067642f
C896 variable_delay_unit_5.tristate_inverter_1.en.n1 VSS 0.85898f
C897 variable_delay_unit_5.tristate_inverter_1.en.n2 VSS 0.944443f
C898 variable_delay_unit_5.tristate_inverter_1.en.t2 VSS 0.093268f
C899 variable_delay_unit_5.tristate_inverter_1.en.t5 VSS 0.086397f
C900 variable_delay_unit_5.tristate_inverter_1.en.t7 VSS 0.093582f
C901 variable_delay_unit_5.tristate_inverter_1.en.n3 VSS 0.091588f
C902 variable_delay_unit_5.tristate_inverter_1.en.n4 VSS 0.06359f
.ends

