magic
tech sky130A
magscale 1 2
timestamp 1729603013
<< error_p >>
rect -29 681 29 687
rect -29 647 -17 681
rect -29 641 29 647
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect -29 -687 29 -681
<< nwell >>
rect -211 -819 211 819
<< pmos >>
rect -15 -600 15 600
<< pdiff >>
rect -73 588 -15 600
rect -73 -588 -61 588
rect -27 -588 -15 588
rect -73 -600 -15 -588
rect 15 588 73 600
rect 15 -588 27 588
rect 61 -588 73 588
rect 15 -600 73 -588
<< pdiffc >>
rect -61 -588 -27 588
rect 27 -588 61 588
<< nsubdiff >>
rect -175 749 -79 783
rect 79 749 175 783
rect -175 687 -141 749
rect 141 687 175 749
rect -175 -749 -141 -687
rect 141 -749 175 -687
rect -175 -783 -79 -749
rect 79 -783 175 -749
<< nsubdiffcont >>
rect -79 749 79 783
rect -175 -687 -141 687
rect 141 -687 175 687
rect -79 -783 79 -749
<< poly >>
rect -33 681 33 697
rect -33 647 -17 681
rect 17 647 33 681
rect -33 631 33 647
rect -15 600 15 631
rect -15 -631 15 -600
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
<< polycont >>
rect -17 647 17 681
rect -17 -681 17 -647
<< locali >>
rect -175 749 -79 783
rect 79 749 175 783
rect -175 687 -141 749
rect 141 687 175 749
rect -33 647 -17 681
rect 17 647 33 681
rect -61 588 -27 604
rect -61 -604 -27 -588
rect 27 588 61 604
rect 27 -604 61 -588
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -175 -749 -141 -687
rect 141 -749 175 -687
rect -175 -783 -79 -749
rect 79 -783 175 -749
<< viali >>
rect -17 647 17 681
rect -61 -588 -27 588
rect 27 -588 61 588
rect -17 -681 17 -647
<< metal1 >>
rect -29 681 29 687
rect -29 647 -17 681
rect 17 647 29 681
rect -29 641 29 647
rect -67 588 -21 600
rect -67 -588 -61 588
rect -27 -588 -21 588
rect -67 -600 -21 -588
rect 21 588 67 600
rect 21 -588 27 588
rect 61 -588 67 588
rect 21 -600 67 -588
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
<< properties >>
string FIXED_BBOX -158 -766 158 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
