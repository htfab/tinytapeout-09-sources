*SWTCH_TWOINV_SKY130NM/SWTCH_TWOINV
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SWTCH_TWOINV_lpe.spi
#else
.include ../../../work/xsch/SWTCH_TWOINV.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VGND  VGND  GND   dc 0
VPWR  VPWR  GND   pwl 0 0 100p {AVDD}

VIN IN GND pwl 0 0 1n 0 2n {AVDD} 3n {AVDD} 4n 0 5n 0 7n {AVDD} 8n {AVDD} 10n 0 

R1 Q_P GND 100k
R2 Q_N GND 100k

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VPWR VGND IN Q_P Q_N SWTCH_TWOINV

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.probe v(VPWR) v(VGND) v(IN) v(Q_P) v(Q_N)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 10n 1p
write
quit
#endif

.endc

.end
