magic
tech sky130A
magscale 1 2
timestamp 1730928108
<< error_p >>
rect -221 522 -163 528
rect -29 522 29 528
rect 163 522 221 528
rect -221 488 -209 522
rect -29 488 -17 522
rect 163 488 175 522
rect -221 482 -163 488
rect -29 482 29 488
rect 163 482 221 488
rect -317 -488 -259 -482
rect -125 -488 -67 -482
rect 67 -488 125 -482
rect 259 -488 317 -482
rect -317 -522 -305 -488
rect -125 -522 -113 -488
rect 67 -522 79 -488
rect 259 -522 271 -488
rect -317 -528 -259 -522
rect -125 -528 -67 -522
rect 67 -528 125 -522
rect 259 -528 317 -522
<< pwell >>
rect -503 -660 503 660
<< nmoslvt >>
rect -303 -450 -273 450
rect -207 -450 -177 450
rect -111 -450 -81 450
rect -15 -450 15 450
rect 81 -450 111 450
rect 177 -450 207 450
rect 273 -450 303 450
<< ndiff >>
rect -365 438 -303 450
rect -365 -438 -353 438
rect -319 -438 -303 438
rect -365 -450 -303 -438
rect -273 438 -207 450
rect -273 -438 -257 438
rect -223 -438 -207 438
rect -273 -450 -207 -438
rect -177 438 -111 450
rect -177 -438 -161 438
rect -127 -438 -111 438
rect -177 -450 -111 -438
rect -81 438 -15 450
rect -81 -438 -65 438
rect -31 -438 -15 438
rect -81 -450 -15 -438
rect 15 438 81 450
rect 15 -438 31 438
rect 65 -438 81 438
rect 15 -450 81 -438
rect 111 438 177 450
rect 111 -438 127 438
rect 161 -438 177 438
rect 111 -450 177 -438
rect 207 438 273 450
rect 207 -438 223 438
rect 257 -438 273 438
rect 207 -450 273 -438
rect 303 438 365 450
rect 303 -438 319 438
rect 353 -438 365 438
rect 303 -450 365 -438
<< ndiffc >>
rect -353 -438 -319 438
rect -257 -438 -223 438
rect -161 -438 -127 438
rect -65 -438 -31 438
rect 31 -438 65 438
rect 127 -438 161 438
rect 223 -438 257 438
rect 319 -438 353 438
<< psubdiff >>
rect -467 590 -371 624
rect 371 590 467 624
rect -467 528 -433 590
rect 433 528 467 590
rect -467 -590 -433 -528
rect 433 -590 467 -528
rect -467 -624 -371 -590
rect 371 -624 467 -590
<< psubdiffcont >>
rect -371 590 371 624
rect -467 -528 -433 528
rect 433 -528 467 528
rect -371 -624 371 -590
<< poly >>
rect -225 522 -159 538
rect -225 488 -209 522
rect -175 488 -159 522
rect -303 450 -273 476
rect -225 472 -159 488
rect -33 522 33 538
rect -33 488 -17 522
rect 17 488 33 522
rect -207 450 -177 472
rect -111 450 -81 476
rect -33 472 33 488
rect 159 522 225 538
rect 159 488 175 522
rect 209 488 225 522
rect -15 450 15 472
rect 81 450 111 476
rect 159 472 225 488
rect 177 450 207 472
rect 273 450 303 476
rect -303 -472 -273 -450
rect -321 -488 -255 -472
rect -207 -476 -177 -450
rect -111 -472 -81 -450
rect -321 -522 -305 -488
rect -271 -522 -255 -488
rect -321 -538 -255 -522
rect -129 -488 -63 -472
rect -15 -476 15 -450
rect 81 -472 111 -450
rect -129 -522 -113 -488
rect -79 -522 -63 -488
rect -129 -538 -63 -522
rect 63 -488 129 -472
rect 177 -476 207 -450
rect 273 -472 303 -450
rect 63 -522 79 -488
rect 113 -522 129 -488
rect 63 -538 129 -522
rect 255 -488 321 -472
rect 255 -522 271 -488
rect 305 -522 321 -488
rect 255 -538 321 -522
<< polycont >>
rect -209 488 -175 522
rect -17 488 17 522
rect 175 488 209 522
rect -305 -522 -271 -488
rect -113 -522 -79 -488
rect 79 -522 113 -488
rect 271 -522 305 -488
<< locali >>
rect -467 590 -371 624
rect 371 590 467 624
rect -467 528 -433 590
rect 433 528 467 590
rect -225 488 -209 522
rect -175 488 -159 522
rect -33 488 -17 522
rect 17 488 33 522
rect 159 488 175 522
rect 209 488 225 522
rect -353 438 -319 454
rect -353 -454 -319 -438
rect -257 438 -223 454
rect -257 -454 -223 -438
rect -161 438 -127 454
rect -161 -454 -127 -438
rect -65 438 -31 454
rect -65 -454 -31 -438
rect 31 438 65 454
rect 31 -454 65 -438
rect 127 438 161 454
rect 127 -454 161 -438
rect 223 438 257 454
rect 223 -454 257 -438
rect 319 438 353 454
rect 319 -454 353 -438
rect -321 -522 -305 -488
rect -271 -522 -255 -488
rect -129 -522 -113 -488
rect -79 -522 -63 -488
rect 63 -522 79 -488
rect 113 -522 129 -488
rect 255 -522 271 -488
rect 305 -522 321 -488
rect -467 -590 -433 -528
rect 433 -590 467 -528
rect -467 -624 -371 -590
rect 371 -624 467 -590
<< viali >>
rect -209 488 -175 522
rect -17 488 17 522
rect 175 488 209 522
rect -353 -438 -319 438
rect -257 -438 -223 438
rect -161 -438 -127 438
rect -65 -438 -31 438
rect 31 -438 65 438
rect 127 -438 161 438
rect 223 -438 257 438
rect 319 -438 353 438
rect -305 -522 -271 -488
rect -113 -522 -79 -488
rect 79 -522 113 -488
rect 271 -522 305 -488
<< metal1 >>
rect -221 522 -163 528
rect -221 488 -209 522
rect -175 488 -163 522
rect -221 482 -163 488
rect -29 522 29 528
rect -29 488 -17 522
rect 17 488 29 522
rect -29 482 29 488
rect 163 522 221 528
rect 163 488 175 522
rect 209 488 221 522
rect 163 482 221 488
rect -359 438 -313 450
rect -359 -438 -353 438
rect -319 -438 -313 438
rect -359 -450 -313 -438
rect -263 438 -217 450
rect -263 -438 -257 438
rect -223 -438 -217 438
rect -263 -450 -217 -438
rect -167 438 -121 450
rect -167 -438 -161 438
rect -127 -438 -121 438
rect -167 -450 -121 -438
rect -71 438 -25 450
rect -71 -438 -65 438
rect -31 -438 -25 438
rect -71 -450 -25 -438
rect 25 438 71 450
rect 25 -438 31 438
rect 65 -438 71 438
rect 25 -450 71 -438
rect 121 438 167 450
rect 121 -438 127 438
rect 161 -438 167 438
rect 121 -450 167 -438
rect 217 438 263 450
rect 217 -438 223 438
rect 257 -438 263 438
rect 217 -450 263 -438
rect 313 438 359 450
rect 313 -438 319 438
rect 353 -438 359 438
rect 313 -450 359 -438
rect -317 -488 -259 -482
rect -317 -522 -305 -488
rect -271 -522 -259 -488
rect -317 -528 -259 -522
rect -125 -488 -67 -482
rect -125 -522 -113 -488
rect -79 -522 -67 -488
rect -125 -528 -67 -522
rect 67 -488 125 -482
rect 67 -522 79 -488
rect 113 -522 125 -488
rect 67 -528 125 -522
rect 259 -488 317 -482
rect 259 -522 271 -488
rect 305 -522 317 -488
rect 259 -528 317 -522
<< properties >>
string FIXED_BBOX -450 -607 450 607
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.5 l 0.150 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
