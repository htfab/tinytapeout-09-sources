magic
tech sky130A
timestamp 1730753331
<< metal1 >>
rect 0 596 27 623
rect 1172 225 1213 227
rect 0 198 53 225
rect 133 198 198 225
rect 278 198 343 225
rect 423 198 488 225
rect 568 198 633 225
rect 713 198 778 225
rect 858 198 923 225
rect 1003 198 1068 225
rect 1148 198 1175 225
rect 1210 198 1213 225
rect 1172 196 1213 198
rect 1317 225 1358 227
rect 1317 198 1320 225
rect 1355 198 1358 225
rect 1317 196 1358 198
rect 1462 225 1503 227
rect 1462 198 1465 225
rect 1500 198 1503 225
rect 1462 196 1503 198
rect 1607 225 1648 227
rect 1607 198 1610 225
rect 1645 198 1648 225
rect 1607 196 1648 198
rect 1728 225 1793 227
rect 1728 198 1755 225
rect 1790 198 1793 225
rect 1728 196 1793 198
rect 1897 225 1938 227
rect 1897 198 1900 225
rect 1935 198 1938 225
rect 1897 196 1938 198
rect 2042 225 2083 227
rect 2042 198 2045 225
rect 2080 198 2083 225
rect 2042 196 2083 198
rect 2187 225 2228 227
rect 2187 198 2190 225
rect 2225 198 2228 225
rect 2187 196 2228 198
rect 2332 225 2373 227
rect 2332 198 2335 225
rect 2370 198 2373 225
rect 2332 196 2373 198
rect 2477 225 2518 227
rect 2477 198 2480 225
rect 2515 198 2518 225
rect 2477 196 2518 198
rect 2622 225 2663 227
rect 2622 198 2625 225
rect 2660 198 2663 225
rect 2622 196 2663 198
rect 2767 225 2808 227
rect 2767 198 2770 225
rect 2805 198 2808 225
rect 2767 196 2808 198
rect 2912 225 2953 227
rect 2912 198 2915 225
rect 2950 198 2953 225
rect 2912 196 2953 198
rect 3057 225 3098 227
rect 3057 198 3060 225
rect 3095 198 3098 225
rect 3057 196 3098 198
rect 3202 225 3243 227
rect 3202 198 3205 225
rect 3240 198 3243 225
rect 3202 196 3243 198
rect 3347 225 3388 227
rect 3347 198 3350 225
rect 3385 198 3388 225
rect 3347 196 3388 198
rect 3492 225 3533 227
rect 3492 198 3495 225
rect 3530 198 3533 225
rect 3492 196 3533 198
rect 3637 225 3678 227
rect 3637 198 3640 225
rect 3675 198 3678 225
rect 3637 196 3678 198
rect 3782 225 3823 227
rect 3782 198 3785 225
rect 3820 198 3823 225
rect 3782 196 3823 198
rect 3927 225 3968 227
rect 3927 198 3930 225
rect 3965 198 3968 225
rect 4025 198 4114 225
rect 3927 196 3968 198
rect 1270 111 1305 114
rect 1270 82 1273 111
rect 1302 82 1305 111
rect 1270 79 1305 82
rect 1415 111 1450 114
rect 1415 82 1418 111
rect 1447 82 1450 111
rect 1415 79 1450 82
rect 1560 111 1595 114
rect 1560 82 1563 111
rect 1592 82 1595 111
rect 1560 79 1595 82
rect 1705 111 1740 114
rect 1705 82 1708 111
rect 1737 82 1740 111
rect 1705 79 1740 82
rect 1850 111 1885 114
rect 1850 82 1853 111
rect 1882 82 1885 111
rect 1850 79 1885 82
rect 1995 111 2030 114
rect 1995 82 1998 111
rect 2027 82 2030 111
rect 1995 79 2030 82
rect 2140 111 2175 114
rect 2140 82 2143 111
rect 2172 82 2175 111
rect 2140 79 2175 82
rect 2285 111 2320 114
rect 2285 82 2288 111
rect 2317 82 2320 111
rect 2285 79 2320 82
rect 2430 111 2465 114
rect 2430 82 2433 111
rect 2462 82 2465 111
rect 2430 79 2465 82
rect 2575 111 2610 114
rect 2575 82 2578 111
rect 2607 82 2610 111
rect 2575 79 2610 82
rect 2720 111 2755 114
rect 2720 82 2723 111
rect 2752 82 2755 111
rect 2720 79 2755 82
rect 2865 111 2900 114
rect 2865 82 2868 111
rect 2897 82 2900 111
rect 2865 79 2900 82
rect 3010 111 3045 114
rect 3010 82 3013 111
rect 3042 82 3045 111
rect 3010 79 3045 82
rect 3155 111 3190 114
rect 3155 82 3158 111
rect 3187 82 3190 111
rect 3155 79 3190 82
rect 3300 111 3335 114
rect 3300 82 3303 111
rect 3332 82 3335 111
rect 3300 79 3335 82
rect 3445 111 3480 114
rect 3445 82 3448 111
rect 3477 82 3480 111
rect 3445 79 3480 82
rect 3590 111 3625 114
rect 3590 82 3593 111
rect 3622 82 3625 111
rect 3590 79 3625 82
rect 3735 111 3770 114
rect 3735 82 3738 111
rect 3767 82 3770 111
rect 3735 79 3770 82
rect 3880 111 3915 114
rect 3880 82 3883 111
rect 3912 82 3915 111
rect 3880 79 3915 82
rect 4025 111 4060 114
rect 4025 82 4028 111
rect 4057 82 4060 111
rect 4025 79 4060 82
rect 0 21 27 48
<< via1 >>
rect 1175 198 1210 225
rect 1320 198 1355 225
rect 1465 198 1500 225
rect 1610 198 1645 225
rect 1755 198 1790 225
rect 1900 198 1935 225
rect 2045 198 2080 225
rect 2190 198 2225 225
rect 2335 198 2370 225
rect 2480 198 2515 225
rect 2625 198 2660 225
rect 2770 198 2805 225
rect 2915 198 2950 225
rect 3060 198 3095 225
rect 3205 198 3240 225
rect 3350 198 3385 225
rect 3495 198 3530 225
rect 3640 198 3675 225
rect 3785 198 3820 225
rect 3930 198 3965 225
rect 1273 82 1302 111
rect 1418 82 1447 111
rect 1563 82 1592 111
rect 1708 82 1737 111
rect 1853 82 1882 111
rect 1998 82 2027 111
rect 2143 82 2172 111
rect 2288 82 2317 111
rect 2433 82 2462 111
rect 2578 82 2607 111
rect 2723 82 2752 111
rect 2868 82 2897 111
rect 3013 82 3042 111
rect 3158 82 3187 111
rect 3303 82 3332 111
rect 3448 82 3477 111
rect 3593 82 3622 111
rect 3738 82 3767 111
rect 3883 82 3912 111
rect 4028 82 4057 111
<< metal2 >>
rect 1172 225 1648 227
rect 1172 198 1175 225
rect 1210 198 1320 225
rect 1355 198 1465 225
rect 1500 198 1610 225
rect 1645 198 1648 225
rect 1172 196 1648 198
rect 1752 225 3968 227
rect 1752 198 1755 225
rect 1790 198 1900 225
rect 1935 198 2045 225
rect 2080 198 2190 225
rect 2225 198 2335 225
rect 2370 198 2480 225
rect 2515 198 2625 225
rect 2660 198 2770 225
rect 2805 198 2915 225
rect 2950 198 3060 225
rect 3095 198 3205 225
rect 3240 198 3350 225
rect 3385 198 3495 225
rect 3530 198 3640 225
rect 3675 198 3785 225
rect 3820 198 3930 225
rect 3965 198 3968 225
rect 1752 196 3968 198
rect 1270 111 1740 114
rect 1270 82 1273 111
rect 1302 82 1418 111
rect 1447 82 1563 111
rect 1592 82 1708 111
rect 1737 82 1740 111
rect 1270 79 1740 82
rect 1850 111 4060 114
rect 1850 82 1853 111
rect 1882 82 1998 111
rect 2027 82 2143 111
rect 2172 82 2288 111
rect 2317 82 2433 111
rect 2462 82 2578 111
rect 2607 82 2723 111
rect 2752 82 2868 111
rect 2897 82 3013 111
rect 3042 82 3158 111
rect 3187 82 3303 111
rect 3332 82 3448 111
rect 3477 82 3593 111
rect 3622 82 3738 111
rect 3767 82 3883 111
rect 3912 82 4028 111
rect 4057 82 4060 111
rect 1850 79 4060 82
use inverter_3_1x4  inverter_3_1x4_0
timestamp 1730750158
transform 1 0 3463 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_1
timestamp 1730750158
transform 1 0 -17 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_2
timestamp 1730750158
transform 1 0 563 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_3
timestamp 1730750158
transform 1 0 1143 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_4
timestamp 1730750158
transform 1 0 1723 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_5
timestamp 1730750158
transform 1 0 2303 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_6
timestamp 1730750158
transform 1 0 2883 0 1 -12
box 17 12 651 653
<< labels >>
rlabel metal1 0 198 27 225 0 stop
port 1 nsew
rlabel metal1 4087 198 4114 225 0 stop_strong
port 2 nsew
rlabel metal1 0 596 27 623 0 VDD
port 3 nsew
rlabel metal1 0 21 27 48 0 VSS
port 4 nsew
<< end >>
