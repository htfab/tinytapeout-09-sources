magic
tech sky130A
timestamp 1731245751
<< metal1 >>
rect 26 779 55 808
rect 73 52 102 81
rect 8841 52 8876 322
<< via1 >>
rect 7493 718 7520 779
<< metal2 >>
rect 161 961 190 990
rect 1640 961 1669 990
rect 3133 961 3162 990
rect 4590 961 4619 990
rect 6044 961 6073 990
rect 58 504 87 533
rect 0 259 29 288
use variable_delay_unit  variable_delay_unit_0
timestamp 1731143787
transform 1 0 700 0 1 52
box -703 -52 850 938
use variable_delay_unit  variable_delay_unit_1
timestamp 1731143787
transform 1 0 2174 0 1 52
box -703 -52 850 938
use variable_delay_unit  variable_delay_unit_2
timestamp 1731143787
transform 1 0 3648 0 1 52
box -703 -52 850 938
use variable_delay_unit  variable_delay_unit_3
timestamp 1731143787
transform 1 0 5122 0 1 52
box -703 -52 850 938
use variable_delay_unit  variable_delay_unit_4
timestamp 1731143787
transform 1 0 6596 0 1 52
box -703 -52 850 938
use variable_delay_unit  variable_delay_unit_5
timestamp 1731143787
transform 1 0 8070 0 1 52
box -703 -52 850 938
<< labels >>
rlabel metal2 58 504 87 533 0 in
port 1 nsew
rlabel metal2 161 961 190 990 0 en_0
port 2 nsew
rlabel metal2 1640 961 1669 990 0 en_1
port 3 nsew
rlabel metal2 3133 961 3162 990 0 en_2
port 4 nsew
rlabel metal2 4590 961 4619 990 0 en_3
port 5 nsew
rlabel metal2 6044 961 6073 990 0 en_4
port 6 nsew
rlabel metal2 0 259 29 288 0 out
port 10 nsew
rlabel metal1 26 779 55 808 0 VDD
port 11 nsew
rlabel metal1 73 52 102 81 0 VSS
port 12 nsew
<< end >>
