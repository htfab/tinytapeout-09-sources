** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/diff_gen.sch
.subckt diff_gen in_delay in_buff out_pos out_neg VDD VSS
*.PININFO VDD:B VSS:B in_delay:I out_pos:O in_buff:I out_neg:O
x1 out_1_1 in_buff in_delay VDD out_2_1 VSS delay_unit
x2 out_1_2 out_1_1 out_2_1 VDD out_2_2 VSS delay_unit
x3 out_1_3 out_1_2 out_2_2 VDD out_2_3 VSS delay_unit
x4 out_1_4 out_1_3 out_2_3 VDD out_2_4 VSS delay_unit
x5 out_1_5 out_1_4 out_2_4 VDD out_2_5 VSS delay_unit
x6 out_1_6 out_1_5 out_2_5 VDD out_2_6 VSS delay_unit
x7 out_pos out_1_6 out_2_6 VDD out_neg VSS delay_unit
.ends

* expanding   symbol:  delay_unit.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/delay_unit.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/delay_unit.sch
.subckt delay_unit out_1 in_1 in_2 VDD out_2 VSS
*.PININFO VDD:B in_1:I out_1:O VSS:B in_2:I out_2:O
XM5 out_2 in_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM7 out_2 in_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM1 out_1 in_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM2 out_1 in_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
XM3 in_1 in_2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM4 in_1 in_2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 in_2 in_1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM8 in_2 in_1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
