* NGSPICE file created from input_stage_parax.ext - technology: sky130A

.subckt input_stage_parax in en t0 t1 t2 t3 VDD VSS out
X0 a_2134_616# t0.t0 a_1870_1170# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X1 a_3160_1170# fine_delay_unit_1.in VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X2 a_3248_1170# fine_delay_unit_1.in a_3160_1170# VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X3 VSS.t13 t3.t0 a_3512_616# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X4 VSS.t21 fine_delay_unit_0.in a_2134_616# VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X5 nand_gate_0.out in.t0 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X6 VSS.t4 fine_delay_unit_1.in a_3512_616# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X7 a_306_476# in.t1 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X8 fine_delay_unit_0.in nand_gate_0.out VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X9 a_3160_1170# fine_delay_unit_1.in a_3248_1170# VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X10 a_2134_616# fine_delay_unit_0.in a_1870_1170# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 VSS.t22 t1.t0 a_2134_616# VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X12 out.t0 a_3160_1170# VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X13 a_3512_616# t2.t0 a_3248_1170# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
X14 a_1870_1170# fine_delay_unit_0.in a_1782_1170# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X15 fine_delay_unit_0.in nand_gate_0.out VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X16 a_3512_616# fine_delay_unit_1.in a_3248_1170# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X17 out.t1 a_3160_1170# VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X18 a_3248_1170# fine_delay_unit_1.in a_3160_1170# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X19 a_1782_1170# fine_delay_unit_0.in VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X20 fine_delay_unit_1.in a_1782_1170# VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X21 VDD.t3 en.t0 nand_gate_0.out VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X22 a_1870_1170# fine_delay_unit_0.in a_1782_1170# VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X23 nand_gate_0.out en.t1 a_306_476# VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X24 a_1782_1170# fine_delay_unit_0.in a_1870_1170# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X25 fine_delay_unit_1.in a_1782_1170# VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
R0 t0 t0.t0 577.703
R1 VSS.n32 VSS.n9 13220.9
R2 VSS.n61 VSS.n33 4447.27
R3 VSS.n48 VSS.n35 4447.27
R4 VSS.n64 VSS.n61 3442.57
R5 VSS.n56 VSS.n35 3442.57
R6 VSS.n33 VSS.n6 3165.68
R7 VSS.n48 VSS.n40 3165.68
R8 VSS.n58 VSS.n57 2206.9
R9 VSS.n64 VSS.n8 2206.4
R10 VSS.n56 VSS.n36 2206.4
R11 VSS.n21 VSS.n18 1707.33
R12 VSS.n21 VSS.n17 1707.33
R13 VSS.n31 VSS.t15 1497.65
R14 VSS.n11 VSS.t15 1497.65
R15 VSS.n68 VSS.n8 1438.1
R16 VSS.n52 VSS.n36 1438.1
R17 VSS.n11 VSS.n9 1366.29
R18 VSS.n19 VSS.n9 1178.35
R19 VSS.n32 VSS.n31 1157.75
R20 VSS.n68 VSS.n6 1065.44
R21 VSS.n52 VSS.n40 1065.44
R22 VSS.n12 VSS.n10 1058.19
R23 VSS.n30 VSS.n10 1058.19
R24 VSS.n65 VSS.n32 1020.69
R25 VSS.t6 VSS.n18 1000.06
R26 VSS.t8 VSS.n19 902.564
R27 VSS.t9 VSS.n48 559.691
R28 VSS.t11 VSS.n58 520.691
R29 VSS.n57 VSS.n34 403.449
R30 VSS.n66 VSS.n65 403.449
R31 VSS.t3 VSS.t9 303.449
R32 VSS.t1 VSS.t3 303.449
R33 VSS.t2 VSS.t5 303.449
R34 VSS.t20 VSS.t11 303.449
R35 VSS.t14 VSS.t20 303.449
R36 VSS.t18 VSS.t17 303.449
R37 VSS.n54 VSS.n36 292.5
R38 VSS.n36 VSS.n34 292.5
R39 VSS.n8 VSS.n7 292.5
R40 VSS.n66 VSS.n8 292.5
R41 VSS.n62 VSS.n5 288.961
R42 VSS.n47 VSS.n37 288.961
R43 VSS.n51 VSS.t0 286.207
R44 VSS.n67 VSS.t19 286.207
R45 VSS.n20 VSS.t8 275.784
R46 VSS.n20 VSS.t6 275.784
R47 VSS.n63 VSS.n62 223.68
R48 VSS.n55 VSS.n37 223.68
R49 VSS.n70 VSS.n5 205.69
R50 VSS.n47 VSS.n39 205.69
R51 VSS.n30 VSS.n29 195
R52 VSS.n31 VSS.n30 195
R53 VSS.n13 VSS.n12 195
R54 VSS.n12 VSS.n11 195
R55 VSS.n49 VSS.t1 155.173
R56 VSS.n60 VSS.t14 155.173
R57 VSS.n53 VSS.n52 146.25
R58 VSS.n52 VSS.n51 146.25
R59 VSS.n69 VSS.n68 146.25
R60 VSS.n68 VSS.n67 146.25
R61 VSS.n28 VSS.n10 146.25
R62 VSS.n10 VSS.t15 146.25
R63 VSS.n63 VSS.n7 143.361
R64 VSS.n55 VSS.n54 143.361
R65 VSS.n22 VSS.n16 110.933
R66 VSS.n22 VSS.n14 110.933
R67 VSS.t0 VSS.n34 103.448
R68 VSS.t19 VSS.n66 103.448
R69 VSS.n17 VSS.n14 97.5005
R70 VSS.n19 VSS.n17 97.5005
R71 VSS.n18 VSS.n16 97.5005
R72 VSS.n69 VSS.n7 93.4405
R73 VSS.n54 VSS.n53 93.4405
R74 VSS.t5 VSS.n50 93.1039
R75 VSS.n59 VSS.t18 93.1039
R76 VSS.n26 VSS.t16 84.1574
R77 VSS.n70 VSS.n69 69.2272
R78 VSS.n53 VSS.n39 69.2272
R79 VSS.n29 VSS.n28 68.7561
R80 VSS.n28 VSS.n13 68.7561
R81 VSS.n42 VSS.n41 67.5509
R82 VSS.n3 VSS.n2 67.5509
R83 VSS.n56 VSS.n55 65.0005
R84 VSS.n57 VSS.n56 65.0005
R85 VSS.n37 VSS.n35 65.0005
R86 VSS.n49 VSS.n35 65.0005
R87 VSS.n64 VSS.n63 65.0005
R88 VSS.n65 VSS.n64 65.0005
R89 VSS.n62 VSS.n61 65.0005
R90 VSS.n61 VSS.n60 65.0005
R91 VSS.n22 VSS.n21 58.5005
R92 VSS.n21 VSS.n20 58.5005
R93 VSS.n50 VSS.n49 55.1729
R94 VSS.n60 VSS.n59 55.1729
R95 VSS.n15 VSS.t7 42.0841
R96 VSS.n42 VSS.t13 41.3938
R97 VSS.n3 VSS.t22 41.3938
R98 VSS.n48 VSS.n47 39.0005
R99 VSS.n33 VSS.n5 39.0005
R100 VSS.n58 VSS.n33 39.0005
R101 VSS.n40 VSS.n39 24.3755
R102 VSS.n50 VSS.n40 24.3755
R103 VSS.n70 VSS.n6 24.3755
R104 VSS.n59 VSS.n6 24.3755
R105 VSS.n41 VSS.t10 17.4005
R106 VSS.n41 VSS.t4 17.4005
R107 VSS.n2 VSS.t12 17.4005
R108 VSS.n2 VSS.t21 17.4005
R109 VSS.n51 VSS.t2 17.2419
R110 VSS.n67 VSS.t17 17.2419
R111 VSS.n29 VSS.n0 3.46248
R112 VSS.n25 VSS.n13 3.46248
R113 VSS.n63 VSS.n1 2.913
R114 VSS.n55 VSS.n38 2.913
R115 VSS.n69 VSS.n1 2.3255
R116 VSS.n53 VSS.n38 2.3255
R117 VSS.n28 VSS.n27 2.3255
R118 VSS.n16 VSS.n15 2.27599
R119 VSS.n24 VSS.n14 2.1305
R120 VSS.n47 VSS.n46 2.12011
R121 VSS.n43 VSS.n5 1.95084
R122 VSS.n23 VSS.n22 1.8605
R123 VSS.n46 VSS.n42 0.957022
R124 VSS.n4 VSS.n3 0.957022
R125 VSS VSS.n0 0.523938
R126 VSS.n25 VSS 0.463123
R127 VSS.n72 VSS.n1 0.440404
R128 VSS.n44 VSS.n38 0.440404
R129 VSS.n45 VSS.n39 0.423227
R130 VSS.n71 VSS.n70 0.423227
R131 VSS.n44 VSS 0.306056
R132 VSS VSS.n72 0.306056
R133 VSS.n24 VSS.n23 0.230892
R134 VSS.n27 VSS.n0 0.189302
R135 VSS.n43 VSS.n4 0.169771
R136 VSS.n46 VSS.n45 0.168035
R137 VSS.n71 VSS.n4 0.168035
R138 VSS VSS.n43 0.15675
R139 VSS.n26 VSS.n25 0.13201
R140 VSS.n23 VSS.n15 0.108343
R141 VSS.n45 VSS.n44 0.104667
R142 VSS.n72 VSS.n71 0.104667
R143 VSS.n27 VSS.n26 0.0577917
R144 VSS VSS.n24 0.0164314
R145 VDD.n45 VDD.n44 1348.04
R146 VDD.n47 VDD.n44 1348.04
R147 VDD.n37 VDD.n35 1307.92
R148 VDD.n23 VDD.n3 1271.17
R149 VDD.n10 VDD.n7 1271.17
R150 VDD.n25 VDD.n3 408.981
R151 VDD.n12 VDD.n7 408.981
R152 VDD.n15 VDD.n14 313.632
R153 VDD.n28 VDD.n27 312.635
R154 VDD.n37 VDD.t10 181.478
R155 VDD.t2 VDD.n45 181.043
R156 VDD.n47 VDD.t8 176.736
R157 VDD.n36 VDD.n33 175.123
R158 VDD.n49 VDD.n48 143.792
R159 VDD.n49 VDD.n42 143.792
R160 VDD.n39 VDD.n33 139.512
R161 VDD.n39 VDD.n38 139.512
R162 VDD.n22 VDD.n2 135.591
R163 VDD.n9 VDD.n6 135.591
R164 VDD.n29 VDD.n0 129.013
R165 VDD.n16 VDD.n4 129.013
R166 VDD.n34 VDD.t11 84.7934
R167 VDD.n43 VDD.t9 84.7879
R168 VDD.n51 VDD.t3 84.7879
R169 VDD.n20 VDD.t7 84.7771
R170 VDD.n8 VDD.t5 84.7771
R171 VDD.n31 VDD.t13 84.7716
R172 VDD.n18 VDD.t1 84.7716
R173 VDD.n28 VDD.n3 61.6672
R174 VDD.n15 VDD.n7 61.6672
R175 VDD.t8 VDD.n46 49.547
R176 VDD.n39 VDD.n35 46.2505
R177 VDD.n46 VDD.t2 45.2386
R178 VDD.n24 VDD.n2 43.625
R179 VDD.n11 VDD.n6 43.625
R180 VDD.n36 VDD.n35 39.3924
R181 VDD.n27 VDD.n0 35.5442
R182 VDD.n14 VDD.n4 35.5275
R183 VDD.n13 VDD.t0 20.8338
R184 VDD.n26 VDD.t12 20.7429
R185 VDD.n38 VDD.n37 20.5561
R186 VDD.n48 VDD.n47 20.5561
R187 VDD.n45 VDD.n42 20.5561
R188 VDD.n25 VDD.n24 20.5561
R189 VDD.n26 VDD.n25 20.5561
R190 VDD.n23 VDD.n22 20.5561
R191 VDD.n26 VDD.n23 20.5561
R192 VDD.n12 VDD.n11 20.5561
R193 VDD.n13 VDD.n12 20.5561
R194 VDD.n10 VDD.n9 20.5561
R195 VDD.n13 VDD.n10 20.5561
R196 VDD.n49 VDD.n44 18.5005
R197 VDD.n46 VDD.n44 18.5005
R198 VDD.n29 VDD.n28 7.70883
R199 VDD.n16 VDD.n15 7.70883
R200 VDD.n29 VDD.n2 6.57828
R201 VDD.n16 VDD.n6 6.57828
R202 VDD.t10 VDD.n36 5.4667
R203 VDD.n14 VDD.n13 5.33119
R204 VDD.n27 VDD.n26 5.31424
R205 VDD.n40 VDD.n39 2.3255
R206 VDD.n41 VDD.n33 2.2281
R207 VDD.n38 VDD.n34 2.17472
R208 VDD.n48 VDD.n43 2.16438
R209 VDD.n9 VDD.n8 2.13168
R210 VDD.t0 VDD.t4 2.08383
R211 VDD.t12 VDD.t6 2.07474
R212 VDD.n52 VDD.n42 2.0406
R213 VDD.n32 VDD.n0 1.96588
R214 VDD.n22 VDD.n21 1.96588
R215 VDD.n19 VDD.n4 1.96588
R216 VDD.n50 VDD.n49 1.8605
R217 VDD.n24 VDD.n1 1.54255
R218 VDD.n11 VDD.n5 1.54255
R219 VDD.n54 VDD.n53 0.6555
R220 VDD.n53 VDD 0.620598
R221 VDD VDD.n54 0.472722
R222 VDD.n21 VDD 0.453625
R223 VDD.n17 VDD.n16 0.423227
R224 VDD.n30 VDD.n29 0.423227
R225 VDD.n53 VDD.n41 0.223
R226 VDD VDD.n19 0.182792
R227 VDD VDD.n32 0.182792
R228 VDD.n21 VDD.n20 0.166299
R229 VDD.n52 VDD.n51 0.129176
R230 VDD.n18 VDD.n17 0.127236
R231 VDD.n31 VDD.n30 0.127236
R232 VDD.n8 VDD.n5 0.115083
R233 VDD.n20 VDD.n1 0.115083
R234 VDD.n50 VDD.n43 0.110794
R235 VDD.n51 VDD.n50 0.105892
R236 VDD.n19 VDD.n18 0.0899097
R237 VDD.n32 VDD.n31 0.0899097
R238 VDD.n17 VDD.n5 0.0647361
R239 VDD.n30 VDD.n1 0.0647361
R240 VDD.n40 VDD.n34 0.0577917
R241 VDD.n54 VDD 0.0439028
R242 VDD VDD.n52 0.0103039
R243 VDD.n41 VDD.n40 0.00440625
R244 t3 t3.t0 727.149
R245 in.n0 in.t0 618.668
R246 in.n0 in.t1 456.997
R247 in in.n0 161.375
R248 t1 t1.t0 727.149
R249 out out.t1 84.8477
R250 out out.t0 84.7009
R251 t2 t2.t0 577.703
R252 en.n0 en.t0 564.04
R253 en.n0 en.t1 511.623
R254 en en.n0 161.333
C0 a_3160_1170# a_3512_616# 0.019821f
C1 a_2134_616# a_1782_1170# 0.019821f
C2 a_1870_1170# t1 0.001628f
C3 t0 t1 0.014805f
C4 a_1870_1170# fine_delay_unit_1.in 7.4e-19
C5 VDD fine_delay_unit_0.in 1.54235f
C6 fine_delay_unit_1.in out 0.00207f
C7 a_2134_616# t2 6.6e-22
C8 nand_gate_0.out fine_delay_unit_0.in 0.062526f
C9 t3 t2 0.014805f
C10 a_1870_1170# en 5.43e-20
C11 a_1782_1170# a_3248_1170# 2.1e-21
C12 t3 a_3248_1170# 0.001628f
C13 t1 a_3512_616# 2.21e-20
C14 t0 a_1870_1170# 0.022005f
C15 t1 fine_delay_unit_0.in 0.020557f
C16 fine_delay_unit_1.in a_3512_616# 0.028846f
C17 fine_delay_unit_1.in fine_delay_unit_0.in 0.030121f
C18 a_3248_1170# t2 0.022005f
C19 a_1782_1170# a_3160_1170# 0.001737f
C20 t3 a_3160_1170# 0.010812f
C21 en fine_delay_unit_0.in 0.001628f
C22 a_1782_1170# VDD 1.25441f
C23 t3 VDD 0.004852f
C24 a_2134_616# nand_gate_0.out 4.47e-20
C25 a_1870_1170# fine_delay_unit_0.in 0.244525f
C26 a_1782_1170# nand_gate_0.out 3.78e-19
C27 out a_3512_616# 7.3e-20
C28 a_3160_1170# t2 0.003337f
C29 t0 fine_delay_unit_0.in 0.009343f
C30 t2 VDD 4.29e-19
C31 a_3248_1170# a_3160_1170# 0.53267f
C32 a_2134_616# t1 0.013742f
C33 a_1782_1170# t1 0.010812f
C34 t1 t3 0.001296f
C35 in VDD 0.118135f
C36 a_2134_616# fine_delay_unit_1.in 5.97e-19
C37 in a_306_476# 0.009499f
C38 a_1782_1170# fine_delay_unit_1.in 0.130035f
C39 in nand_gate_0.out 0.050326f
C40 fine_delay_unit_1.in t3 0.020481f
C41 t1 t2 5.63e-19
C42 fine_delay_unit_1.in t2 0.009158f
C43 a_3160_1170# VDD 1.25072f
C44 a_2134_616# a_1870_1170# 0.556904f
C45 t1 a_3248_1170# 1.01e-19
C46 a_1870_1170# a_1782_1170# 0.53267f
C47 t0 a_2134_616# 0.02185f
C48 t0 a_1782_1170# 0.003337f
C49 out t3 0.034216f
C50 fine_delay_unit_1.in a_3248_1170# 0.244525f
C51 VDD a_306_476# 7.57e-19
C52 nand_gate_0.out VDD 1.28298f
C53 nand_gate_0.out a_306_476# 0.355469f
C54 t0 t2 0.003859f
C55 in en 0.078266f
C56 fine_delay_unit_1.in a_3160_1170# 0.253736f
C57 a_1782_1170# a_3512_616# 7.57e-22
C58 a_2134_616# fine_delay_unit_0.in 0.028846f
C59 out a_3248_1170# 3.44e-20
C60 t3 a_3512_616# 0.013742f
C61 a_1782_1170# fine_delay_unit_0.in 0.253714f
C62 t1 VDD 0.003164f
C63 nand_gate_0.out t1 2.7e-20
C64 fine_delay_unit_1.in VDD 1.33558f
C65 t2 a_3512_616# 0.02185f
C66 out a_3160_1170# 0.115353f
C67 en VDD 0.150039f
C68 en a_306_476# 0.009499f
C69 nand_gate_0.out en 0.12418f
C70 a_3248_1170# a_3512_616# 0.556904f
C71 a_3248_1170# fine_delay_unit_0.in 1.39e-20
C72 in fine_delay_unit_0.in 5.53e-19
C73 t0 VDD 6.26e-19
C74 fine_delay_unit_1.in t1 0.039118f
C75 a_1870_1170# nand_gate_0.out 5.26e-20
C76 out VDD 0.963042f
C77 t0 nand_gate_0.out 9.64e-20
C78 t2 VSS 0.309129f
C79 t3 VSS 0.375997f
C80 t0 VSS 0.309038f
C81 t1 VSS 0.371058f
C82 out VSS 0.493979f
C83 en VSS 0.179937f
C84 in VSS 0.247895f
C85 VDD VSS 11.680599f
C86 a_3512_616# VSS 0.612975f
C87 a_3248_1170# VSS 0.387205f
C88 a_2134_616# VSS 0.612975f
C89 a_1870_1170# VSS 0.387205f
C90 a_306_476# VSS 0.371906f
C91 a_3160_1170# VSS 0.739963f
C92 fine_delay_unit_1.in VSS 1.71608f
C93 nand_gate_0.out VSS 0.89651f
C94 a_1782_1170# VSS 0.7316f
C95 fine_delay_unit_0.in VSS 1.83203f
.ends

