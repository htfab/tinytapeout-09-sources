magic
tech sky130A
timestamp 1730835638
<< metal1 >>
rect 0 605 18 623
rect 157 225 198 227
rect 0 198 53 225
rect 133 198 160 225
rect 195 198 198 225
rect 157 196 198 198
rect 302 225 343 227
rect 302 198 305 225
rect 340 198 343 225
rect 302 196 343 198
rect 447 225 488 227
rect 447 198 450 225
rect 485 198 488 225
rect 447 196 488 198
rect 592 225 633 227
rect 737 225 778 227
rect 592 198 595 225
rect 630 198 633 225
rect 713 198 740 225
rect 775 198 778 225
rect 592 196 633 198
rect 737 196 778 198
rect 882 225 923 227
rect 882 198 885 225
rect 920 198 923 225
rect 882 196 923 198
rect 1027 225 1068 227
rect 1027 198 1030 225
rect 1065 198 1068 225
rect 1148 198 1214 225
rect 1027 196 1068 198
rect 255 111 290 114
rect 255 82 258 111
rect 287 82 290 111
rect 255 79 290 82
rect 400 111 435 114
rect 400 82 403 111
rect 432 82 435 111
rect 400 79 435 82
rect 545 111 580 114
rect 545 82 548 111
rect 577 82 580 111
rect 545 79 580 82
rect 690 111 725 114
rect 690 82 693 111
rect 722 82 725 111
rect 690 79 725 82
rect 835 111 870 114
rect 835 82 838 111
rect 867 82 870 111
rect 835 79 870 82
rect 980 111 1015 114
rect 980 82 983 111
rect 1012 82 1015 111
rect 980 79 1015 82
rect 1125 111 1160 114
rect 1125 82 1128 111
rect 1157 82 1160 111
rect 1125 79 1160 82
rect 0 30 18 48
<< via1 >>
rect 160 198 195 225
rect 305 198 340 225
rect 450 198 485 225
rect 595 198 630 225
rect 740 198 775 225
rect 885 198 920 225
rect 1030 198 1065 225
rect 258 82 287 111
rect 403 82 432 111
rect 548 82 577 111
rect 693 82 722 111
rect 838 82 867 111
rect 983 82 1012 111
rect 1128 82 1157 111
<< metal2 >>
rect 157 225 633 227
rect 157 198 160 225
rect 195 198 305 225
rect 340 198 450 225
rect 485 198 595 225
rect 630 198 633 225
rect 157 196 633 198
rect 737 225 1068 227
rect 737 198 740 225
rect 775 198 885 225
rect 920 198 1030 225
rect 1065 198 1068 225
rect 737 196 1068 198
rect 255 111 725 114
rect 255 82 258 111
rect 287 82 403 111
rect 432 82 548 111
rect 577 82 693 111
rect 722 82 725 111
rect 255 79 725 82
rect 835 111 1160 114
rect 835 82 838 111
rect 867 82 983 111
rect 1012 82 1128 111
rect 1157 82 1160 111
rect 835 79 1160 82
use inverter_3_1x4  inverter_3_1x4_0
timestamp 1730750158
transform 1 0 -17 0 1 -12
box 17 12 651 653
use inverter_3_1x4  inverter_3_1x4_1
timestamp 1730750158
transform 1 0 563 0 1 -12
box 17 12 651 653
<< labels >>
rlabel metal1 0 198 27 225 0 start
port 1 nsew
rlabel metal1 1187 198 1214 225 0 start_delay
port 2 nsew
rlabel metal2 690 79 725 114 0 start_buff
port 3 nsew
rlabel metal1 0 605 18 623 0 VDD
port 4 nsew
rlabel metal1 0 30 18 48 0 VSS
port 5 nsew
<< end >>
