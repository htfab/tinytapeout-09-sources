magic
tech sky130A
magscale 1 2
timestamp 1730308116
<< error_p >>
rect -1031 34 -961 36
rect -865 34 -795 36
rect -699 34 -629 36
rect -533 34 -463 36
rect -367 34 -297 36
rect -201 34 -131 36
rect -35 34 35 36
rect 131 34 201 36
rect 297 34 367 36
rect 463 34 533 36
rect 629 34 699 36
rect 795 34 865 36
rect 961 34 1031 36
<< pwell >>
rect -1197 -632 1197 632
<< psubdiff >>
rect -1161 562 -1065 596
rect 1065 562 1161 596
rect -1161 500 -1127 562
rect 1127 500 1161 562
rect -1161 -562 -1127 -500
rect 1127 -562 1161 -500
rect -1161 -596 -1065 -562
rect 1065 -596 1161 -562
<< psubdiffcont >>
rect -1065 562 1065 596
rect -1161 -500 -1127 500
rect 1127 -500 1161 500
rect -1065 -596 1065 -562
<< xpolycontact >>
rect -1031 34 -961 466
rect -1031 -466 -961 -34
rect -865 34 -795 466
rect -865 -466 -795 -34
rect -699 34 -629 466
rect -699 -466 -629 -34
rect -533 34 -463 466
rect -533 -466 -463 -34
rect -367 34 -297 466
rect -367 -466 -297 -34
rect -201 34 -131 466
rect -201 -466 -131 -34
rect -35 34 35 466
rect -35 -466 35 -34
rect 131 34 201 466
rect 131 -466 201 -34
rect 297 34 367 466
rect 297 -466 367 -34
rect 463 34 533 466
rect 463 -466 533 -34
rect 629 34 699 466
rect 629 -466 699 -34
rect 795 34 865 466
rect 795 -466 865 -34
rect 961 34 1031 466
rect 961 -466 1031 -34
<< xpolyres >>
rect -1031 -34 -961 34
rect -865 -34 -795 34
rect -699 -34 -629 34
rect -533 -34 -463 34
rect -367 -34 -297 34
rect -201 -34 -131 34
rect -35 -34 35 34
rect 131 -34 201 34
rect 297 -34 367 34
rect 463 -34 533 34
rect 629 -34 699 34
rect 795 -34 865 34
rect 961 -34 1031 34
<< locali >>
rect -1161 562 -1065 596
rect 1065 562 1161 596
rect -1161 500 -1127 562
rect 1127 500 1161 562
rect -1161 -562 -1127 -500
rect 1127 -562 1161 -500
rect -1161 -596 -1065 -562
rect 1065 -596 1161 -562
<< viali >>
rect -1015 51 -977 448
rect -849 51 -811 448
rect -683 51 -645 448
rect -517 51 -479 448
rect -351 51 -313 448
rect -185 51 -147 448
rect -19 51 19 448
rect 147 51 185 448
rect 313 51 351 448
rect 479 51 517 448
rect 645 51 683 448
rect 811 51 849 448
rect 977 51 1015 448
rect -1015 -448 -977 -51
rect -849 -448 -811 -51
rect -683 -448 -645 -51
rect -517 -448 -479 -51
rect -351 -448 -313 -51
rect -185 -448 -147 -51
rect -19 -448 19 -51
rect 147 -448 185 -51
rect 313 -448 351 -51
rect 479 -448 517 -51
rect 645 -448 683 -51
rect 811 -448 849 -51
rect 977 -448 1015 -51
<< metal1 >>
rect -1021 448 -971 460
rect -1021 51 -1015 448
rect -977 51 -971 448
rect -1021 39 -971 51
rect -855 448 -805 460
rect -855 51 -849 448
rect -811 51 -805 448
rect -855 39 -805 51
rect -689 448 -639 460
rect -689 51 -683 448
rect -645 51 -639 448
rect -689 39 -639 51
rect -523 448 -473 460
rect -523 51 -517 448
rect -479 51 -473 448
rect -523 39 -473 51
rect -357 448 -307 460
rect -357 51 -351 448
rect -313 51 -307 448
rect -357 39 -307 51
rect -191 448 -141 460
rect -191 51 -185 448
rect -147 51 -141 448
rect -191 39 -141 51
rect -25 448 25 460
rect -25 51 -19 448
rect 19 51 25 448
rect -25 39 25 51
rect 141 448 191 460
rect 141 51 147 448
rect 185 51 191 448
rect 141 39 191 51
rect 307 448 357 460
rect 307 51 313 448
rect 351 51 357 448
rect 307 39 357 51
rect 473 448 523 460
rect 473 51 479 448
rect 517 51 523 448
rect 473 39 523 51
rect 639 448 689 460
rect 639 51 645 448
rect 683 51 689 448
rect 639 39 689 51
rect 805 448 855 460
rect 805 51 811 448
rect 849 51 855 448
rect 805 39 855 51
rect 971 448 1021 460
rect 971 51 977 448
rect 1015 51 1021 448
rect 971 39 1021 51
rect -1021 -51 -971 -39
rect -1021 -448 -1015 -51
rect -977 -448 -971 -51
rect -1021 -460 -971 -448
rect -855 -51 -805 -39
rect -855 -448 -849 -51
rect -811 -448 -805 -51
rect -855 -460 -805 -448
rect -689 -51 -639 -39
rect -689 -448 -683 -51
rect -645 -448 -639 -51
rect -689 -460 -639 -448
rect -523 -51 -473 -39
rect -523 -448 -517 -51
rect -479 -448 -473 -51
rect -523 -460 -473 -448
rect -357 -51 -307 -39
rect -357 -448 -351 -51
rect -313 -448 -307 -51
rect -357 -460 -307 -448
rect -191 -51 -141 -39
rect -191 -448 -185 -51
rect -147 -448 -141 -51
rect -191 -460 -141 -448
rect -25 -51 25 -39
rect -25 -448 -19 -51
rect 19 -448 25 -51
rect -25 -460 25 -448
rect 141 -51 191 -39
rect 141 -448 147 -51
rect 185 -448 191 -51
rect 141 -460 191 -448
rect 307 -51 357 -39
rect 307 -448 313 -51
rect 351 -448 357 -51
rect 307 -460 357 -448
rect 473 -51 523 -39
rect 473 -448 479 -51
rect 517 -448 523 -51
rect 473 -460 523 -448
rect 639 -51 689 -39
rect 639 -448 645 -51
rect 683 -448 689 -51
rect 639 -460 689 -448
rect 805 -51 855 -39
rect 805 -448 811 -51
rect 849 -448 855 -51
rect 805 -460 855 -448
rect 971 -51 1021 -39
rect 971 -448 977 -51
rect 1015 -448 1021 -51
rect 971 -460 1021 -448
<< properties >>
string FIXED_BBOX -1144 -579 1144 579
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.50 m 1 nx 13 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
