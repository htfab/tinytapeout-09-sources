** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/fine_delay.sch
.subckt fine_delay in t0 t1 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B t0:I t1:I
XM1 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net3 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net3 t1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM8 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM9 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net2 in net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net2 t0 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
