magic
tech sky130A
magscale 1 2
timestamp 1730892491
<< nwell >>
rect -996 -419 996 419
<< pmos >>
rect -800 -200 800 200
<< pdiff >>
rect -858 188 -800 200
rect -858 -188 -846 188
rect -812 -188 -800 188
rect -858 -200 -800 -188
rect 800 188 858 200
rect 800 -188 812 188
rect 846 -188 858 188
rect 800 -200 858 -188
<< pdiffc >>
rect -846 -188 -812 188
rect 812 -188 846 188
<< nsubdiff >>
rect -960 349 -864 383
rect 864 349 960 383
rect -960 287 -926 349
rect 926 287 960 349
rect -960 -349 -926 -287
rect 926 -349 960 -287
rect -960 -383 -864 -349
rect 864 -383 960 -349
<< nsubdiffcont >>
rect -864 349 864 383
rect -960 -287 -926 287
rect 926 -287 960 287
rect -864 -383 864 -349
<< poly >>
rect -800 281 800 297
rect -800 247 -784 281
rect 784 247 800 281
rect -800 200 800 247
rect -800 -247 800 -200
rect -800 -281 -784 -247
rect 784 -281 800 -247
rect -800 -297 800 -281
<< polycont >>
rect -784 247 784 281
rect -784 -281 784 -247
<< locali >>
rect -960 349 -864 383
rect 864 349 960 383
rect -960 287 -926 349
rect 926 287 960 349
rect -800 247 -784 281
rect 784 247 800 281
rect -846 188 -812 204
rect -846 -204 -812 -188
rect 812 188 846 204
rect 812 -204 846 -188
rect -800 -281 -784 -247
rect 784 -281 800 -247
rect -960 -349 -926 -287
rect 926 -349 960 -287
rect -960 -383 -864 -349
rect 864 -383 960 -349
<< viali >>
rect -784 247 784 281
rect -846 -188 -812 188
rect 812 -188 846 188
rect -784 -281 784 -247
<< metal1 >>
rect -796 281 796 287
rect -796 247 -784 281
rect 784 247 796 281
rect -796 241 796 247
rect -852 188 -806 200
rect -852 -188 -846 188
rect -812 -188 -806 188
rect -852 -200 -806 -188
rect 806 188 852 200
rect 806 -188 812 188
rect 846 -188 852 188
rect 806 -200 852 -188
rect -796 -247 796 -241
rect -796 -281 -784 -247
rect 784 -281 796 -247
rect -796 -287 796 -281
<< properties >>
string FIXED_BBOX -943 -366 943 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 8.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
