** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_short.sch
.subckt variable_delay_short in en_0 en_1 en_2 en_3 en_4 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en_0:I en_1:I en_2:I en_3:I en_4:I
x1 in en_0 out_1 forward_0 out VDD VSS variable_delay_unit
x2 forward_0 en_1 out_2 forward_1 out_1 VDD VSS variable_delay_unit
x3 forward_1 en_2 out_3 forward_2 out_2 VDD VSS variable_delay_unit
x4 forward_2 en_3 out_4 forward_3 out_3 VDD VSS variable_delay_unit
x9 forward_4 VDD VSS net1 out_5 VDD VSS variable_delay_unit
x5 forward_3 en_4 out_5 forward_4 out_4 VDD VSS variable_delay_unit
.ends

* expanding   symbol:  variable_delay_unit.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_unit.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/variable_delay_unit.sch
.subckt variable_delay_unit in en back forward out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en:I back:I forward:O
x1 forward en nen out VDD VSS tristate_inverter
x2 in forward VDD VSS inverter_2
x3 en nen VDD VSS inverter_2
x4 back nen en out VDD VSS tristate_inverter
.ends


* expanding   symbol:  tristate_inverter.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tristate_inverter.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/tristate_inverter.sch
.subckt tristate_inverter in en nen out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B en:I nen:I
XM5 out in net2 VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM7 out in net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 net2 nen VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=9 nf=1 m=1
XM2 net1 en VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=3 nf=1 m=1
.ends


* expanding   symbol:  inverter_2.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sch
.subckt inverter_2 in out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
