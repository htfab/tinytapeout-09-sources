VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt09ball4_logo
  CLASS BLOCK ;
  FOREIGN tt09ball4_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 92.400 BY 29.400 ;
  OBS
      LAYER met1 ;
        RECT 0.000 28.840 92.400 29.400 ;
        RECT 0.000 28.560 44.240 28.840 ;
      LAYER met1 ;
        RECT 44.240 28.560 45.080 28.840 ;
      LAYER met1 ;
        RECT 45.080 28.560 92.400 28.840 ;
        RECT 0.000 26.040 43.960 28.560 ;
      LAYER met1 ;
        RECT 43.960 28.280 45.920 28.560 ;
      LAYER met1 ;
        RECT 45.920 28.280 92.400 28.560 ;
      LAYER met1 ;
        RECT 43.960 26.040 44.520 28.280 ;
      LAYER met1 ;
        RECT 44.520 28.000 45.080 28.280 ;
      LAYER met1 ;
        RECT 45.080 28.000 46.480 28.280 ;
      LAYER met1 ;
        RECT 46.480 28.000 92.400 28.280 ;
        RECT 44.520 27.720 45.920 28.000 ;
      LAYER met1 ;
        RECT 45.920 27.720 47.320 28.000 ;
      LAYER met1 ;
        RECT 47.320 27.720 92.400 28.000 ;
        RECT 44.520 27.440 46.480 27.720 ;
      LAYER met1 ;
        RECT 46.480 27.440 47.880 27.720 ;
      LAYER met1 ;
        RECT 47.880 27.440 53.760 27.720 ;
      LAYER met1 ;
        RECT 53.760 27.440 56.280 27.720 ;
      LAYER met1 ;
        RECT 56.280 27.440 92.400 27.720 ;
        RECT 44.520 27.160 47.320 27.440 ;
      LAYER met1 ;
        RECT 47.320 27.160 48.440 27.440 ;
      LAYER met1 ;
        RECT 48.440 27.160 52.360 27.440 ;
      LAYER met1 ;
        RECT 52.360 27.160 56.560 27.440 ;
      LAYER met1 ;
        RECT 44.520 26.880 47.880 27.160 ;
      LAYER met1 ;
        RECT 47.880 26.880 49.000 27.160 ;
      LAYER met1 ;
        RECT 49.000 26.880 49.280 27.160 ;
      LAYER met1 ;
        RECT 49.280 26.880 50.400 27.160 ;
      LAYER met1 ;
        RECT 50.400 26.880 51.240 27.160 ;
      LAYER met1 ;
        RECT 51.240 26.880 53.760 27.160 ;
      LAYER met1 ;
        RECT 53.760 26.880 56.000 27.160 ;
        RECT 44.520 26.600 48.440 26.880 ;
      LAYER met1 ;
        RECT 48.440 26.600 52.360 26.880 ;
      LAYER met1 ;
        RECT 52.360 26.600 56.000 26.880 ;
        RECT 44.520 26.320 48.720 26.600 ;
      LAYER met1 ;
        RECT 48.720 26.320 49.560 26.600 ;
      LAYER met1 ;
        RECT 49.560 26.320 50.120 26.600 ;
      LAYER met1 ;
        RECT 50.120 26.320 51.240 26.600 ;
      LAYER met1 ;
        RECT 51.240 26.320 56.000 26.600 ;
        RECT 44.520 26.040 48.440 26.320 ;
      LAYER met1 ;
        RECT 48.440 26.040 50.960 26.320 ;
      LAYER met1 ;
        RECT 50.960 26.040 56.000 26.320 ;
        RECT 0.000 25.760 43.400 26.040 ;
      LAYER met1 ;
        RECT 43.400 25.760 44.520 26.040 ;
      LAYER met1 ;
        RECT 44.520 25.760 47.040 26.040 ;
      LAYER met1 ;
        RECT 47.040 25.760 52.080 26.040 ;
      LAYER met1 ;
        RECT 52.080 25.760 56.000 26.040 ;
        RECT 0.000 25.480 42.840 25.760 ;
      LAYER met1 ;
        RECT 42.840 25.480 43.960 25.760 ;
      LAYER met1 ;
        RECT 43.960 25.480 44.240 25.760 ;
        RECT 0.000 25.200 5.880 25.480 ;
      LAYER met1 ;
        RECT 5.880 25.200 9.800 25.480 ;
      LAYER met1 ;
        RECT 9.800 25.200 23.240 25.480 ;
      LAYER met1 ;
        RECT 23.240 25.200 27.160 25.480 ;
      LAYER met1 ;
        RECT 27.160 25.200 42.280 25.480 ;
      LAYER met1 ;
        RECT 42.280 25.200 43.400 25.480 ;
      LAYER met1 ;
        RECT 43.400 25.200 44.240 25.480 ;
      LAYER met1 ;
        RECT 44.240 25.200 44.800 25.760 ;
      LAYER met1 ;
        RECT 44.800 25.480 45.920 25.760 ;
      LAYER met1 ;
        RECT 45.920 25.480 48.440 25.760 ;
      LAYER met1 ;
        RECT 48.440 25.480 50.960 25.760 ;
      LAYER met1 ;
        RECT 50.960 25.480 52.640 25.760 ;
      LAYER met1 ;
        RECT 52.640 25.480 56.000 25.760 ;
        RECT 44.800 25.200 45.080 25.480 ;
      LAYER met1 ;
        RECT 45.080 25.200 47.040 25.480 ;
      LAYER met1 ;
        RECT 47.040 25.200 52.080 25.480 ;
      LAYER met1 ;
        RECT 52.080 25.200 53.200 25.480 ;
      LAYER met1 ;
        RECT 53.200 25.200 56.000 25.480 ;
      LAYER met1 ;
        RECT 56.000 25.200 56.560 27.160 ;
      LAYER met1 ;
        RECT 56.560 25.200 92.400 27.440 ;
        RECT 0.000 24.920 5.040 25.200 ;
      LAYER met1 ;
        RECT 5.040 24.920 10.360 25.200 ;
      LAYER met1 ;
        RECT 10.360 24.920 22.400 25.200 ;
      LAYER met1 ;
        RECT 22.400 24.920 28.000 25.200 ;
      LAYER met1 ;
        RECT 28.000 24.920 42.000 25.200 ;
      LAYER met1 ;
        RECT 42.000 24.920 42.840 25.200 ;
      LAYER met1 ;
        RECT 42.840 24.920 44.240 25.200 ;
      LAYER met1 ;
        RECT 44.240 24.920 45.920 25.200 ;
      LAYER met1 ;
        RECT 45.920 24.920 52.640 25.200 ;
      LAYER met1 ;
        RECT 52.640 24.920 53.760 25.200 ;
      LAYER met1 ;
        RECT 53.760 24.920 55.720 25.200 ;
        RECT 0.000 24.640 4.480 24.920 ;
      LAYER met1 ;
        RECT 4.480 24.640 10.920 24.920 ;
      LAYER met1 ;
        RECT 10.920 24.640 21.840 24.920 ;
      LAYER met1 ;
        RECT 21.840 24.640 28.560 24.920 ;
      LAYER met1 ;
        RECT 28.560 24.640 41.720 24.920 ;
      LAYER met1 ;
        RECT 41.720 24.640 42.560 24.920 ;
      LAYER met1 ;
        RECT 42.560 24.640 43.960 24.920 ;
      LAYER met1 ;
        RECT 43.960 24.640 45.080 24.920 ;
      LAYER met1 ;
        RECT 45.080 24.640 53.200 24.920 ;
      LAYER met1 ;
        RECT 53.200 24.640 54.040 24.920 ;
      LAYER met1 ;
        RECT 54.040 24.640 55.720 24.920 ;
      LAYER met1 ;
        RECT 55.720 24.640 56.280 25.200 ;
      LAYER met1 ;
        RECT 56.280 24.640 92.400 25.200 ;
        RECT 0.000 24.360 3.920 24.640 ;
      LAYER met1 ;
        RECT 3.920 24.360 11.480 24.640 ;
      LAYER met1 ;
        RECT 11.480 24.360 21.280 24.640 ;
      LAYER met1 ;
        RECT 21.280 24.360 29.120 24.640 ;
      LAYER met1 ;
        RECT 29.120 24.360 41.720 24.640 ;
      LAYER met1 ;
        RECT 41.720 24.360 43.120 24.640 ;
      LAYER met1 ;
        RECT 43.120 24.360 43.680 24.640 ;
      LAYER met1 ;
        RECT 43.680 24.360 44.520 24.640 ;
      LAYER met1 ;
        RECT 44.520 24.360 53.480 24.640 ;
      LAYER met1 ;
        RECT 53.480 24.360 54.320 24.640 ;
      LAYER met1 ;
        RECT 54.320 24.360 55.440 24.640 ;
      LAYER met1 ;
        RECT 55.440 24.360 56.560 24.640 ;
      LAYER met1 ;
        RECT 56.560 24.360 92.400 24.640 ;
        RECT 0.000 24.080 3.360 24.360 ;
      LAYER met1 ;
        RECT 3.360 24.080 6.160 24.360 ;
      LAYER met1 ;
        RECT 6.160 24.080 9.240 24.360 ;
      LAYER met1 ;
        RECT 9.240 24.080 12.040 24.360 ;
      LAYER met1 ;
        RECT 12.040 24.080 21.000 24.360 ;
      LAYER met1 ;
        RECT 21.000 24.080 23.800 24.360 ;
      LAYER met1 ;
        RECT 23.800 24.080 26.600 24.360 ;
      LAYER met1 ;
        RECT 26.600 24.080 29.400 24.360 ;
      LAYER met1 ;
        RECT 29.400 24.080 42.560 24.360 ;
      LAYER met1 ;
        RECT 42.560 24.080 44.240 24.360 ;
      LAYER met1 ;
        RECT 44.240 24.080 54.040 24.360 ;
      LAYER met1 ;
        RECT 54.040 24.080 54.600 24.360 ;
      LAYER met1 ;
        RECT 54.600 24.080 55.440 24.360 ;
      LAYER met1 ;
        RECT 55.440 24.080 56.840 24.360 ;
      LAYER met1 ;
        RECT 56.840 24.080 92.400 24.360 ;
        RECT 0.000 23.800 3.080 24.080 ;
      LAYER met1 ;
        RECT 3.080 23.800 5.320 24.080 ;
      LAYER met1 ;
        RECT 5.320 23.800 10.080 24.080 ;
      LAYER met1 ;
        RECT 10.080 23.800 12.320 24.080 ;
      LAYER met1 ;
        RECT 12.320 23.800 20.720 24.080 ;
      LAYER met1 ;
        RECT 20.720 23.800 22.960 24.080 ;
      LAYER met1 ;
        RECT 22.960 23.800 27.440 24.080 ;
      LAYER met1 ;
        RECT 27.440 23.800 29.680 24.080 ;
      LAYER met1 ;
        RECT 29.680 23.800 42.840 24.080 ;
      LAYER met1 ;
        RECT 42.840 23.800 43.680 24.080 ;
      LAYER met1 ;
        RECT 43.680 23.800 54.320 24.080 ;
      LAYER met1 ;
        RECT 54.320 23.800 54.880 24.080 ;
      LAYER met1 ;
        RECT 54.880 23.800 55.160 24.080 ;
      LAYER met1 ;
        RECT 55.160 23.800 56.000 24.080 ;
      LAYER met1 ;
        RECT 56.000 23.800 56.280 24.080 ;
      LAYER met1 ;
        RECT 56.280 23.800 57.120 24.080 ;
      LAYER met1 ;
        RECT 57.120 23.800 92.400 24.080 ;
        RECT 0.000 23.520 2.800 23.800 ;
      LAYER met1 ;
        RECT 2.800 23.520 4.760 23.800 ;
      LAYER met1 ;
        RECT 4.760 23.520 10.640 23.800 ;
      LAYER met1 ;
        RECT 10.640 23.520 12.600 23.800 ;
      LAYER met1 ;
        RECT 12.600 23.520 20.440 23.800 ;
      LAYER met1 ;
        RECT 20.440 23.520 22.400 23.800 ;
      LAYER met1 ;
        RECT 22.400 23.520 28.000 23.800 ;
      LAYER met1 ;
        RECT 28.000 23.520 29.960 23.800 ;
      LAYER met1 ;
        RECT 29.960 23.520 42.560 23.800 ;
      LAYER met1 ;
        RECT 42.560 23.520 43.400 23.800 ;
      LAYER met1 ;
        RECT 43.400 23.520 54.600 23.800 ;
      LAYER met1 ;
        RECT 54.600 23.520 55.720 23.800 ;
      LAYER met1 ;
        RECT 55.720 23.520 56.560 23.800 ;
      LAYER met1 ;
        RECT 56.560 23.520 57.400 23.800 ;
      LAYER met1 ;
        RECT 57.400 23.520 92.400 23.800 ;
        RECT 0.000 23.240 2.520 23.520 ;
      LAYER met1 ;
        RECT 2.520 23.240 4.480 23.520 ;
      LAYER met1 ;
        RECT 4.480 23.240 10.920 23.520 ;
      LAYER met1 ;
        RECT 10.920 23.240 12.880 23.520 ;
      LAYER met1 ;
        RECT 12.880 23.240 20.160 23.520 ;
      LAYER met1 ;
        RECT 20.160 23.240 21.840 23.520 ;
      LAYER met1 ;
        RECT 21.840 23.240 28.560 23.520 ;
      LAYER met1 ;
        RECT 28.560 23.240 30.240 23.520 ;
      LAYER met1 ;
        RECT 30.240 23.240 42.560 23.520 ;
        RECT 0.000 22.960 2.240 23.240 ;
      LAYER met1 ;
        RECT 2.240 22.960 3.920 23.240 ;
      LAYER met1 ;
        RECT 3.920 22.960 11.480 23.240 ;
      LAYER met1 ;
        RECT 11.480 22.960 13.160 23.240 ;
      LAYER met1 ;
        RECT 13.160 22.960 19.880 23.240 ;
      LAYER met1 ;
        RECT 19.880 22.960 21.560 23.240 ;
      LAYER met1 ;
        RECT 21.560 22.960 28.840 23.240 ;
      LAYER met1 ;
        RECT 28.840 22.960 30.520 23.240 ;
      LAYER met1 ;
        RECT 30.520 22.960 42.560 23.240 ;
      LAYER met1 ;
        RECT 42.560 22.960 43.120 23.520 ;
      LAYER met1 ;
        RECT 43.120 22.960 54.880 23.520 ;
      LAYER met1 ;
        RECT 54.880 22.960 55.440 23.520 ;
      LAYER met1 ;
        RECT 55.440 23.240 56.840 23.520 ;
      LAYER met1 ;
        RECT 56.840 23.240 57.680 23.520 ;
      LAYER met1 ;
        RECT 57.680 23.240 92.400 23.520 ;
        RECT 55.440 22.960 57.120 23.240 ;
      LAYER met1 ;
        RECT 57.120 22.960 57.960 23.240 ;
      LAYER met1 ;
        RECT 57.960 22.960 92.400 23.240 ;
        RECT 0.000 22.680 1.960 22.960 ;
      LAYER met1 ;
        RECT 1.960 22.680 3.640 22.960 ;
      LAYER met1 ;
        RECT 3.640 22.680 11.760 22.960 ;
      LAYER met1 ;
        RECT 11.760 22.680 13.440 22.960 ;
      LAYER met1 ;
        RECT 13.440 22.680 19.600 22.960 ;
      LAYER met1 ;
        RECT 19.600 22.680 21.280 22.960 ;
      LAYER met1 ;
        RECT 21.280 22.680 29.120 22.960 ;
      LAYER met1 ;
        RECT 29.120 22.680 30.800 22.960 ;
      LAYER met1 ;
        RECT 30.800 22.680 42.280 22.960 ;
        RECT 0.000 22.120 1.680 22.680 ;
      LAYER met1 ;
        RECT 1.680 22.120 8.960 22.680 ;
      LAYER met1 ;
        RECT 8.960 22.400 12.040 22.680 ;
      LAYER met1 ;
        RECT 12.040 22.400 13.440 22.680 ;
      LAYER met1 ;
        RECT 13.440 22.400 19.320 22.680 ;
      LAYER met1 ;
        RECT 19.320 22.400 21.000 22.680 ;
      LAYER met1 ;
        RECT 21.000 22.400 24.920 22.680 ;
      LAYER met1 ;
        RECT 24.920 22.400 26.040 22.680 ;
      LAYER met1 ;
        RECT 26.040 22.400 29.400 22.680 ;
      LAYER met1 ;
        RECT 29.400 22.400 31.080 22.680 ;
      LAYER met1 ;
        RECT 31.080 22.400 42.280 22.680 ;
        RECT 0.000 21.560 1.400 22.120 ;
      LAYER met1 ;
        RECT 1.400 21.560 8.960 22.120 ;
      LAYER met1 ;
        RECT 8.960 21.840 12.320 22.400 ;
      LAYER met1 ;
        RECT 12.320 22.120 13.720 22.400 ;
      LAYER met1 ;
        RECT 13.720 22.120 19.320 22.400 ;
      LAYER met1 ;
        RECT 19.320 22.120 20.720 22.400 ;
      LAYER met1 ;
        RECT 20.720 22.120 24.080 22.400 ;
      LAYER met1 ;
        RECT 24.080 22.120 26.880 22.400 ;
      LAYER met1 ;
        RECT 26.880 22.120 29.680 22.400 ;
      LAYER met1 ;
        RECT 29.680 22.120 31.360 22.400 ;
      LAYER met1 ;
        RECT 31.360 22.120 42.280 22.400 ;
      LAYER met1 ;
        RECT 42.280 22.120 42.840 22.960 ;
      LAYER met1 ;
        RECT 42.840 22.680 55.160 22.960 ;
      LAYER met1 ;
        RECT 55.160 22.680 55.720 22.960 ;
      LAYER met1 ;
        RECT 55.720 22.680 57.120 22.960 ;
      LAYER met1 ;
        RECT 57.120 22.680 58.240 22.960 ;
      LAYER met1 ;
        RECT 42.840 22.400 55.440 22.680 ;
        RECT 42.840 22.120 47.040 22.400 ;
      LAYER met1 ;
        RECT 47.040 22.120 47.320 22.400 ;
      LAYER met1 ;
        RECT 47.320 22.120 55.440 22.400 ;
      LAYER met1 ;
        RECT 55.440 22.120 56.000 22.680 ;
      LAYER met1 ;
        RECT 56.000 22.400 56.560 22.680 ;
      LAYER met1 ;
        RECT 56.560 22.400 58.240 22.680 ;
      LAYER met1 ;
        RECT 58.240 22.400 92.400 22.960 ;
        RECT 56.000 22.120 56.280 22.400 ;
      LAYER met1 ;
        RECT 56.280 22.120 57.400 22.400 ;
      LAYER met1 ;
        RECT 57.400 22.120 71.960 22.400 ;
      LAYER met1 ;
        RECT 71.960 22.120 72.800 22.400 ;
      LAYER met1 ;
        RECT 72.800 22.120 92.400 22.400 ;
      LAYER met1 ;
        RECT 12.320 21.840 14.000 22.120 ;
      LAYER met1 ;
        RECT 14.000 21.840 19.040 22.120 ;
      LAYER met1 ;
        RECT 19.040 21.840 20.440 22.120 ;
      LAYER met1 ;
        RECT 20.440 21.840 23.520 22.120 ;
      LAYER met1 ;
        RECT 23.520 21.840 27.160 22.120 ;
      LAYER met1 ;
        RECT 27.160 21.840 29.960 22.120 ;
      LAYER met1 ;
        RECT 29.960 21.840 31.360 22.120 ;
      LAYER met1 ;
        RECT 31.360 21.840 42.000 22.120 ;
      LAYER met1 ;
        RECT 42.000 21.840 42.840 22.120 ;
      LAYER met1 ;
        RECT 42.840 21.840 44.520 22.120 ;
      LAYER met1 ;
        RECT 44.520 21.840 44.800 22.120 ;
      LAYER met1 ;
        RECT 44.800 21.840 45.920 22.120 ;
      LAYER met1 ;
        RECT 45.920 21.840 46.200 22.120 ;
      LAYER met1 ;
        RECT 8.960 21.560 12.600 21.840 ;
      LAYER met1 ;
        RECT 12.600 21.560 14.000 21.840 ;
      LAYER met1 ;
        RECT 14.000 21.560 18.760 21.840 ;
        RECT 0.000 20.720 1.120 21.560 ;
      LAYER met1 ;
        RECT 1.120 20.720 8.960 21.560 ;
      LAYER met1 ;
        RECT 8.960 21.000 12.880 21.560 ;
      LAYER met1 ;
        RECT 12.880 21.000 14.280 21.560 ;
      LAYER met1 ;
        RECT 14.280 21.000 18.760 21.560 ;
      LAYER met1 ;
        RECT 18.760 21.280 20.160 21.840 ;
      LAYER met1 ;
        RECT 20.160 21.560 23.240 21.840 ;
      LAYER met1 ;
        RECT 23.240 21.560 27.440 21.840 ;
      LAYER met1 ;
        RECT 27.440 21.560 30.240 21.840 ;
        RECT 20.160 21.280 22.960 21.560 ;
      LAYER met1 ;
        RECT 22.960 21.280 27.720 21.560 ;
      LAYER met1 ;
        RECT 27.720 21.280 30.240 21.560 ;
      LAYER met1 ;
        RECT 30.240 21.280 31.640 21.840 ;
      LAYER met1 ;
        RECT 31.640 21.560 42.000 21.840 ;
      LAYER met1 ;
        RECT 42.000 21.560 42.560 21.840 ;
      LAYER met1 ;
        RECT 31.640 21.280 41.720 21.560 ;
      LAYER met1 ;
        RECT 41.720 21.280 42.560 21.560 ;
      LAYER met1 ;
        RECT 42.560 21.280 44.240 21.840 ;
      LAYER met1 ;
        RECT 44.240 21.280 44.800 21.840 ;
      LAYER met1 ;
        RECT 44.800 21.560 45.640 21.840 ;
      LAYER met1 ;
        RECT 45.640 21.560 46.200 21.840 ;
      LAYER met1 ;
        RECT 46.200 21.560 46.760 22.120 ;
      LAYER met1 ;
        RECT 46.760 21.560 47.320 22.120 ;
      LAYER met1 ;
        RECT 47.320 21.840 49.280 22.120 ;
      LAYER met1 ;
        RECT 49.280 21.840 49.840 22.120 ;
      LAYER met1 ;
        RECT 49.840 21.840 55.720 22.120 ;
      LAYER met1 ;
        RECT 55.720 21.840 56.840 22.120 ;
      LAYER met1 ;
        RECT 56.840 21.840 71.680 22.120 ;
      LAYER met1 ;
        RECT 71.680 21.840 72.800 22.120 ;
      LAYER met1 ;
        RECT 72.800 21.840 79.520 22.120 ;
      LAYER met1 ;
        RECT 79.520 21.840 80.080 22.120 ;
      LAYER met1 ;
        RECT 80.080 21.840 91.000 22.120 ;
      LAYER met1 ;
        RECT 91.000 21.840 91.560 22.120 ;
      LAYER met1 ;
        RECT 91.560 21.840 92.400 22.120 ;
        RECT 47.320 21.560 49.000 21.840 ;
      LAYER met1 ;
        RECT 49.000 21.560 49.840 21.840 ;
      LAYER met1 ;
        RECT 49.840 21.560 50.680 21.840 ;
      LAYER met1 ;
        RECT 50.680 21.560 50.960 21.840 ;
      LAYER met1 ;
        RECT 50.960 21.560 52.080 21.840 ;
      LAYER met1 ;
        RECT 52.080 21.560 52.360 21.840 ;
      LAYER met1 ;
        RECT 52.360 21.560 55.720 21.840 ;
      LAYER met1 ;
        RECT 18.760 21.000 19.880 21.280 ;
      LAYER met1 ;
        RECT 19.880 21.000 22.960 21.280 ;
      LAYER met1 ;
        RECT 22.960 21.000 28.000 21.280 ;
      LAYER met1 ;
        RECT 8.960 20.720 13.160 21.000 ;
      LAYER met1 ;
        RECT 13.160 20.720 14.280 21.000 ;
      LAYER met1 ;
        RECT 14.280 20.720 18.480 21.000 ;
      LAYER met1 ;
        RECT 18.480 20.720 19.880 21.000 ;
      LAYER met1 ;
        RECT 19.880 20.720 22.680 21.000 ;
      LAYER met1 ;
        RECT 22.680 20.720 24.920 21.000 ;
      LAYER met1 ;
        RECT 24.920 20.720 26.040 21.000 ;
      LAYER met1 ;
        RECT 26.040 20.720 28.000 21.000 ;
      LAYER met1 ;
        RECT 28.000 20.720 30.520 21.280 ;
      LAYER met1 ;
        RECT 30.520 20.720 31.920 21.280 ;
      LAYER met1 ;
        RECT 31.920 21.000 41.720 21.280 ;
      LAYER met1 ;
        RECT 41.720 21.000 42.280 21.280 ;
      LAYER met1 ;
        RECT 31.920 20.720 41.440 21.000 ;
      LAYER met1 ;
        RECT 41.440 20.720 42.280 21.000 ;
      LAYER met1 ;
        RECT 42.280 20.720 43.960 21.280 ;
      LAYER met1 ;
        RECT 43.960 20.720 44.800 21.280 ;
      LAYER met1 ;
        RECT 44.800 21.000 45.360 21.560 ;
      LAYER met1 ;
        RECT 45.360 21.000 46.200 21.560 ;
      LAYER met1 ;
        RECT 46.200 21.000 46.480 21.560 ;
      LAYER met1 ;
        RECT 46.480 21.000 47.600 21.560 ;
      LAYER met1 ;
        RECT 47.600 21.280 48.720 21.560 ;
      LAYER met1 ;
        RECT 48.720 21.280 50.120 21.560 ;
      LAYER met1 ;
        RECT 47.600 21.000 48.440 21.280 ;
      LAYER met1 ;
        RECT 48.440 21.000 49.280 21.280 ;
      LAYER met1 ;
        RECT 49.280 21.000 49.560 21.280 ;
      LAYER met1 ;
        RECT 49.560 21.000 50.120 21.280 ;
      LAYER met1 ;
        RECT 50.120 21.000 50.680 21.560 ;
      LAYER met1 ;
        RECT 50.680 21.280 51.520 21.560 ;
      LAYER met1 ;
        RECT 51.520 21.280 52.080 21.560 ;
      LAYER met1 ;
        RECT 52.080 21.280 52.640 21.560 ;
      LAYER met1 ;
        RECT 52.640 21.280 55.720 21.560 ;
      LAYER met1 ;
        RECT 55.720 21.280 56.560 21.840 ;
      LAYER met1 ;
        RECT 56.560 21.560 70.840 21.840 ;
      LAYER met1 ;
        RECT 70.840 21.560 73.080 21.840 ;
      LAYER met1 ;
        RECT 73.080 21.560 79.520 21.840 ;
      LAYER met1 ;
        RECT 79.520 21.560 80.920 21.840 ;
      LAYER met1 ;
        RECT 80.920 21.560 90.160 21.840 ;
      LAYER met1 ;
        RECT 90.160 21.560 91.840 21.840 ;
      LAYER met1 ;
        RECT 56.560 21.280 70.000 21.560 ;
      LAYER met1 ;
        RECT 70.000 21.280 73.360 21.560 ;
      LAYER met1 ;
        RECT 73.360 21.280 77.560 21.560 ;
      LAYER met1 ;
        RECT 77.560 21.280 78.400 21.560 ;
      LAYER met1 ;
        RECT 78.400 21.280 79.520 21.560 ;
      LAYER met1 ;
        RECT 50.680 21.000 51.800 21.280 ;
      LAYER met1 ;
        RECT 51.800 21.000 52.360 21.280 ;
        RECT 44.800 20.720 45.080 21.000 ;
      LAYER met1 ;
        RECT 45.080 20.720 47.600 21.000 ;
      LAYER met1 ;
        RECT 47.600 20.720 48.160 21.000 ;
      LAYER met1 ;
        RECT 48.160 20.720 49.000 21.000 ;
      LAYER met1 ;
        RECT 49.000 20.720 49.560 21.000 ;
      LAYER met1 ;
        RECT 49.560 20.720 52.080 21.000 ;
      LAYER met1 ;
        RECT 52.080 20.720 52.360 21.000 ;
      LAYER met1 ;
        RECT 52.360 20.720 52.920 21.280 ;
      LAYER met1 ;
        RECT 52.920 21.000 56.000 21.280 ;
      LAYER met1 ;
        RECT 56.000 21.000 56.840 21.280 ;
      LAYER met1 ;
        RECT 56.840 21.000 68.880 21.280 ;
      LAYER met1 ;
        RECT 68.880 21.000 73.080 21.280 ;
      LAYER met1 ;
        RECT 73.080 21.000 77.560 21.280 ;
        RECT 52.920 20.720 56.280 21.000 ;
        RECT 0.000 20.160 4.760 20.720 ;
        RECT 0.000 19.600 0.840 20.160 ;
      LAYER met1 ;
        RECT 0.840 19.600 1.960 20.160 ;
      LAYER met1 ;
        RECT 0.000 17.640 0.560 19.600 ;
      LAYER met1 ;
        RECT 0.560 19.320 1.960 19.600 ;
      LAYER met1 ;
        RECT 1.960 19.320 4.760 20.160 ;
      LAYER met1 ;
        RECT 4.760 19.320 7.000 20.720 ;
      LAYER met1 ;
        RECT 7.000 20.440 13.160 20.720 ;
      LAYER met1 ;
        RECT 13.160 20.440 14.560 20.720 ;
      LAYER met1 ;
        RECT 7.000 19.320 13.440 20.440 ;
      LAYER met1 ;
        RECT 13.440 19.600 14.560 20.440 ;
      LAYER met1 ;
        RECT 14.560 20.160 18.480 20.720 ;
      LAYER met1 ;
        RECT 18.480 20.160 19.600 20.720 ;
      LAYER met1 ;
        RECT 19.600 20.440 22.680 20.720 ;
      LAYER met1 ;
        RECT 22.680 20.440 24.640 20.720 ;
      LAYER met1 ;
        RECT 24.640 20.440 26.320 20.720 ;
        RECT 14.560 19.600 18.200 20.160 ;
      LAYER met1 ;
        RECT 18.200 19.600 19.600 20.160 ;
      LAYER met1 ;
        RECT 19.600 19.600 22.400 20.440 ;
      LAYER met1 ;
        RECT 13.440 19.320 14.840 19.600 ;
        RECT 0.560 17.920 1.680 19.320 ;
      LAYER met1 ;
        RECT 1.680 17.920 4.760 19.320 ;
      LAYER met1 ;
        RECT 0.560 17.640 1.960 17.920 ;
      LAYER met1 ;
        RECT 0.000 16.240 0.840 17.640 ;
      LAYER met1 ;
        RECT 0.840 16.800 1.960 17.640 ;
      LAYER met1 ;
        RECT 1.960 16.800 4.760 17.920 ;
      LAYER met1 ;
        RECT 4.760 17.360 12.320 19.320 ;
      LAYER met1 ;
        RECT 12.320 17.640 13.720 19.320 ;
      LAYER met1 ;
        RECT 13.720 17.640 14.840 19.320 ;
      LAYER met1 ;
        RECT 12.320 17.360 13.440 17.640 ;
      LAYER met1 ;
        RECT 13.440 17.360 14.840 17.640 ;
      LAYER met1 ;
        RECT 14.840 17.360 18.200 19.600 ;
      LAYER met1 ;
        RECT 18.200 17.360 19.320 19.600 ;
      LAYER met1 ;
        RECT 19.320 19.040 22.400 19.600 ;
      LAYER met1 ;
        RECT 22.400 19.320 24.360 20.440 ;
      LAYER met1 ;
        RECT 24.360 19.320 26.320 20.440 ;
      LAYER met1 ;
        RECT 26.320 19.880 28.280 20.720 ;
      LAYER met1 ;
        RECT 28.280 19.880 30.800 20.720 ;
      LAYER met1 ;
        RECT 30.800 20.440 31.920 20.720 ;
      LAYER met1 ;
        RECT 31.920 20.440 41.160 20.720 ;
      LAYER met1 ;
        RECT 41.160 20.440 42.000 20.720 ;
      LAYER met1 ;
        RECT 42.000 20.440 43.680 20.720 ;
      LAYER met1 ;
        RECT 43.680 20.440 46.760 20.720 ;
      LAYER met1 ;
        RECT 46.760 20.440 47.040 20.720 ;
      LAYER met1 ;
        RECT 47.040 20.440 47.600 20.720 ;
      LAYER met1 ;
        RECT 47.600 20.440 47.880 20.720 ;
      LAYER met1 ;
        RECT 47.880 20.440 48.720 20.720 ;
      LAYER met1 ;
        RECT 48.720 20.440 49.560 20.720 ;
      LAYER met1 ;
        RECT 49.560 20.440 50.960 20.720 ;
      LAYER met1 ;
        RECT 50.960 20.440 51.520 20.720 ;
      LAYER met1 ;
        RECT 51.520 20.440 53.200 20.720 ;
      LAYER met1 ;
        RECT 53.200 20.440 54.040 20.720 ;
      LAYER met1 ;
        RECT 54.040 20.440 54.320 20.720 ;
      LAYER met1 ;
        RECT 54.320 20.440 56.280 20.720 ;
      LAYER met1 ;
        RECT 30.800 19.880 32.200 20.440 ;
      LAYER met1 ;
        RECT 32.200 20.160 41.160 20.440 ;
      LAYER met1 ;
        RECT 41.160 20.160 41.720 20.440 ;
      LAYER met1 ;
        RECT 41.720 20.160 43.400 20.440 ;
      LAYER met1 ;
        RECT 43.400 20.160 45.360 20.440 ;
      LAYER met1 ;
        RECT 45.360 20.160 45.640 20.440 ;
      LAYER met1 ;
        RECT 22.400 19.040 24.640 19.320 ;
      LAYER met1 ;
        RECT 24.640 19.040 26.320 19.320 ;
      LAYER met1 ;
        RECT 26.320 19.040 28.560 19.880 ;
      LAYER met1 ;
        RECT 19.320 18.480 22.680 19.040 ;
      LAYER met1 ;
        RECT 22.680 18.760 24.920 19.040 ;
      LAYER met1 ;
        RECT 24.920 18.760 26.040 19.040 ;
      LAYER met1 ;
        RECT 26.040 18.760 28.560 19.040 ;
        RECT 22.680 18.480 28.560 18.760 ;
      LAYER met1 ;
        RECT 19.320 17.920 22.960 18.480 ;
      LAYER met1 ;
        RECT 22.960 18.200 28.560 18.480 ;
      LAYER met1 ;
        RECT 28.560 18.200 31.080 19.880 ;
      LAYER met1 ;
        RECT 22.960 17.920 28.280 18.200 ;
      LAYER met1 ;
        RECT 19.320 17.640 23.240 17.920 ;
      LAYER met1 ;
        RECT 23.240 17.640 28.280 17.920 ;
      LAYER met1 ;
        RECT 19.320 17.360 23.800 17.640 ;
      LAYER met1 ;
        RECT 23.800 17.360 25.760 17.640 ;
      LAYER met1 ;
        RECT 25.760 17.360 26.320 17.640 ;
      LAYER met1 ;
        RECT 26.320 17.360 28.280 17.640 ;
      LAYER met1 ;
        RECT 28.280 17.360 31.080 18.200 ;
      LAYER met1 ;
        RECT 31.080 17.360 32.200 19.880 ;
      LAYER met1 ;
        RECT 32.200 19.040 40.880 20.160 ;
      LAYER met1 ;
        RECT 40.880 19.880 41.720 20.160 ;
      LAYER met1 ;
        RECT 41.720 19.880 43.120 20.160 ;
      LAYER met1 ;
        RECT 43.120 19.880 45.080 20.160 ;
      LAYER met1 ;
        RECT 45.080 19.880 45.640 20.160 ;
      LAYER met1 ;
        RECT 45.640 19.880 46.480 20.440 ;
      LAYER met1 ;
        RECT 46.480 19.880 47.040 20.440 ;
      LAYER met1 ;
        RECT 47.040 20.160 48.440 20.440 ;
      LAYER met1 ;
        RECT 48.440 20.160 49.560 20.440 ;
      LAYER met1 ;
        RECT 49.560 20.160 50.400 20.440 ;
      LAYER met1 ;
        RECT 50.400 20.160 52.080 20.440 ;
      LAYER met1 ;
        RECT 52.080 20.160 53.480 20.440 ;
      LAYER met1 ;
        RECT 53.480 20.160 54.040 20.440 ;
      LAYER met1 ;
        RECT 54.040 20.160 54.600 20.440 ;
      LAYER met1 ;
        RECT 54.600 20.160 56.280 20.440 ;
      LAYER met1 ;
        RECT 56.280 20.160 56.840 21.000 ;
      LAYER met1 ;
        RECT 56.840 20.160 67.760 21.000 ;
      LAYER met1 ;
        RECT 67.760 20.720 72.800 21.000 ;
      LAYER met1 ;
        RECT 72.800 20.720 77.560 21.000 ;
      LAYER met1 ;
        RECT 47.040 19.880 48.160 20.160 ;
      LAYER met1 ;
        RECT 48.160 19.880 52.360 20.160 ;
      LAYER met1 ;
        RECT 52.360 19.880 53.480 20.160 ;
      LAYER met1 ;
        RECT 53.480 19.880 54.320 20.160 ;
      LAYER met1 ;
        RECT 54.320 19.880 54.600 20.160 ;
      LAYER met1 ;
        RECT 54.600 19.880 56.560 20.160 ;
      LAYER met1 ;
        RECT 40.880 19.320 41.440 19.880 ;
      LAYER met1 ;
        RECT 41.440 19.600 42.840 19.880 ;
      LAYER met1 ;
        RECT 42.840 19.600 44.800 19.880 ;
      LAYER met1 ;
        RECT 44.800 19.600 45.640 19.880 ;
      LAYER met1 ;
        RECT 45.640 19.600 46.200 19.880 ;
      LAYER met1 ;
        RECT 46.200 19.600 47.320 19.880 ;
        RECT 41.440 19.320 41.720 19.600 ;
      LAYER met1 ;
        RECT 41.720 19.320 42.280 19.600 ;
      LAYER met1 ;
        RECT 42.280 19.320 42.560 19.600 ;
      LAYER met1 ;
        RECT 42.560 19.320 43.680 19.600 ;
        RECT 40.880 19.040 43.680 19.320 ;
      LAYER met1 ;
        RECT 32.200 18.480 41.160 19.040 ;
      LAYER met1 ;
        RECT 41.160 18.760 42.560 19.040 ;
        RECT 41.160 18.480 41.720 18.760 ;
      LAYER met1 ;
        RECT 41.720 18.480 42.000 18.760 ;
        RECT 32.200 18.200 42.000 18.480 ;
      LAYER met1 ;
        RECT 42.000 18.200 42.560 18.760 ;
      LAYER met1 ;
        RECT 42.560 18.200 42.840 19.040 ;
        RECT 32.200 17.360 41.720 18.200 ;
      LAYER met1 ;
        RECT 41.720 17.360 42.280 18.200 ;
      LAYER met1 ;
        RECT 42.280 17.360 42.840 18.200 ;
      LAYER met1 ;
        RECT 42.840 17.920 43.680 19.040 ;
      LAYER met1 ;
        RECT 43.680 17.920 43.960 19.600 ;
      LAYER met1 ;
        RECT 42.840 17.360 43.400 17.920 ;
        RECT 0.840 16.240 2.240 16.800 ;
      LAYER met1 ;
        RECT 0.000 15.680 1.120 16.240 ;
      LAYER met1 ;
        RECT 1.120 15.960 2.240 16.240 ;
      LAYER met1 ;
        RECT 2.240 15.960 4.760 16.800 ;
      LAYER met1 ;
        RECT 4.760 15.960 7.000 17.360 ;
      LAYER met1 ;
        RECT 7.000 15.960 8.120 17.360 ;
      LAYER met1 ;
        RECT 1.120 15.680 2.520 15.960 ;
      LAYER met1 ;
        RECT 2.520 15.680 8.120 15.960 ;
        RECT 0.000 15.120 1.400 15.680 ;
      LAYER met1 ;
        RECT 1.400 15.120 2.800 15.680 ;
      LAYER met1 ;
        RECT 2.800 15.120 8.120 15.680 ;
        RECT 0.000 14.560 1.680 15.120 ;
      LAYER met1 ;
        RECT 1.680 14.840 3.080 15.120 ;
      LAYER met1 ;
        RECT 3.080 14.840 8.120 15.120 ;
      LAYER met1 ;
        RECT 1.680 14.560 3.360 14.840 ;
      LAYER met1 ;
        RECT 3.360 14.560 8.120 14.840 ;
        RECT 0.000 14.280 1.960 14.560 ;
      LAYER met1 ;
        RECT 1.960 14.280 3.640 14.560 ;
      LAYER met1 ;
        RECT 3.640 14.280 8.120 14.560 ;
        RECT 0.000 14.000 2.240 14.280 ;
      LAYER met1 ;
        RECT 2.240 14.000 3.920 14.280 ;
      LAYER met1 ;
        RECT 3.920 14.000 8.120 14.280 ;
        RECT 0.000 13.720 2.520 14.000 ;
      LAYER met1 ;
        RECT 2.520 13.720 4.200 14.000 ;
      LAYER met1 ;
        RECT 4.200 13.720 8.120 14.000 ;
        RECT 0.000 13.440 2.800 13.720 ;
      LAYER met1 ;
        RECT 2.800 13.440 4.480 13.720 ;
      LAYER met1 ;
        RECT 4.480 13.440 8.120 13.720 ;
        RECT 0.000 13.160 3.080 13.440 ;
      LAYER met1 ;
        RECT 3.080 13.160 5.040 13.440 ;
      LAYER met1 ;
        RECT 5.040 13.160 8.120 13.440 ;
        RECT 0.000 12.880 3.360 13.160 ;
      LAYER met1 ;
        RECT 3.360 12.880 5.600 13.160 ;
      LAYER met1 ;
        RECT 5.600 12.880 8.120 13.160 ;
        RECT 0.000 12.600 3.640 12.880 ;
      LAYER met1 ;
        RECT 3.640 12.600 7.000 12.880 ;
      LAYER met1 ;
        RECT 7.000 12.600 8.120 12.880 ;
      LAYER met1 ;
        RECT 8.120 12.600 10.360 17.360 ;
      LAYER met1 ;
        RECT 10.360 16.800 13.440 17.360 ;
      LAYER met1 ;
        RECT 13.440 16.800 14.560 17.360 ;
      LAYER met1 ;
        RECT 14.560 16.800 18.200 17.360 ;
      LAYER met1 ;
        RECT 18.200 16.800 19.600 17.360 ;
      LAYER met1 ;
        RECT 19.600 17.080 26.320 17.360 ;
      LAYER met1 ;
        RECT 26.320 17.080 28.000 17.360 ;
      LAYER met1 ;
        RECT 19.600 16.800 26.040 17.080 ;
      LAYER met1 ;
        RECT 26.040 16.800 28.000 17.080 ;
      LAYER met1 ;
        RECT 28.000 16.800 30.800 17.360 ;
      LAYER met1 ;
        RECT 30.800 16.800 32.200 17.360 ;
      LAYER met1 ;
        RECT 32.200 16.800 41.440 17.360 ;
      LAYER met1 ;
        RECT 41.440 17.080 42.280 17.360 ;
      LAYER met1 ;
        RECT 42.280 17.080 42.560 17.360 ;
      LAYER met1 ;
        RECT 42.560 17.080 43.400 17.360 ;
      LAYER met1 ;
        RECT 43.400 17.080 43.960 17.920 ;
        RECT 10.360 15.960 13.160 16.800 ;
      LAYER met1 ;
        RECT 13.160 16.240 14.560 16.800 ;
      LAYER met1 ;
        RECT 14.560 16.240 18.480 16.800 ;
      LAYER met1 ;
        RECT 18.480 16.520 19.600 16.800 ;
      LAYER met1 ;
        RECT 19.600 16.520 25.760 16.800 ;
      LAYER met1 ;
        RECT 25.760 16.520 27.720 16.800 ;
        RECT 13.160 15.960 14.280 16.240 ;
      LAYER met1 ;
        RECT 14.280 15.960 18.480 16.240 ;
      LAYER met1 ;
        RECT 18.480 15.960 19.880 16.520 ;
      LAYER met1 ;
        RECT 19.880 16.240 25.200 16.520 ;
      LAYER met1 ;
        RECT 25.200 16.240 27.720 16.520 ;
      LAYER met1 ;
        RECT 27.720 16.240 30.800 16.800 ;
      LAYER met1 ;
        RECT 30.800 16.240 31.920 16.800 ;
      LAYER met1 ;
        RECT 19.880 15.960 24.360 16.240 ;
      LAYER met1 ;
        RECT 24.360 15.960 27.440 16.240 ;
      LAYER met1 ;
        RECT 27.440 15.960 30.520 16.240 ;
      LAYER met1 ;
        RECT 30.520 15.960 31.920 16.240 ;
      LAYER met1 ;
        RECT 31.920 15.960 41.440 16.800 ;
      LAYER met1 ;
        RECT 41.440 15.960 42.000 17.080 ;
      LAYER met1 ;
        RECT 42.000 16.800 42.560 17.080 ;
      LAYER met1 ;
        RECT 42.560 16.800 43.120 17.080 ;
      LAYER met1 ;
        RECT 42.000 15.960 42.280 16.800 ;
      LAYER met1 ;
        RECT 42.280 16.240 43.120 16.800 ;
      LAYER met1 ;
        RECT 43.120 16.240 43.960 17.080 ;
      LAYER met1 ;
        RECT 42.280 15.960 42.840 16.240 ;
      LAYER met1 ;
        RECT 10.360 15.400 12.880 15.960 ;
      LAYER met1 ;
        RECT 12.880 15.680 14.280 15.960 ;
      LAYER met1 ;
        RECT 14.280 15.680 18.760 15.960 ;
      LAYER met1 ;
        RECT 18.760 15.680 19.880 15.960 ;
      LAYER met1 ;
        RECT 19.880 15.680 23.240 15.960 ;
      LAYER met1 ;
        RECT 23.240 15.680 27.160 15.960 ;
      LAYER met1 ;
        RECT 27.160 15.680 30.520 15.960 ;
      LAYER met1 ;
        RECT 30.520 15.680 31.640 15.960 ;
        RECT 12.880 15.400 14.000 15.680 ;
      LAYER met1 ;
        RECT 14.000 15.400 18.760 15.680 ;
      LAYER met1 ;
        RECT 18.760 15.400 20.160 15.680 ;
      LAYER met1 ;
        RECT 20.160 15.400 23.240 15.680 ;
      LAYER met1 ;
        RECT 23.240 15.400 26.880 15.680 ;
      LAYER met1 ;
        RECT 26.880 15.400 30.240 15.680 ;
      LAYER met1 ;
        RECT 30.240 15.400 31.640 15.680 ;
      LAYER met1 ;
        RECT 31.640 15.400 41.440 15.960 ;
      LAYER met1 ;
        RECT 41.440 15.400 42.840 15.960 ;
      LAYER met1 ;
        RECT 42.840 15.400 43.960 16.240 ;
      LAYER met1 ;
        RECT 43.960 15.400 44.520 19.600 ;
      LAYER met1 ;
        RECT 44.520 19.320 47.320 19.600 ;
      LAYER met1 ;
        RECT 47.320 19.320 48.160 19.880 ;
      LAYER met1 ;
        RECT 48.160 19.600 52.640 19.880 ;
      LAYER met1 ;
        RECT 52.640 19.600 53.760 19.880 ;
      LAYER met1 ;
        RECT 53.760 19.600 54.320 19.880 ;
      LAYER met1 ;
        RECT 54.320 19.600 54.880 19.880 ;
      LAYER met1 ;
        RECT 48.160 19.320 52.920 19.600 ;
      LAYER met1 ;
        RECT 52.920 19.320 54.040 19.600 ;
      LAYER met1 ;
        RECT 54.040 19.320 54.600 19.600 ;
        RECT 44.520 18.760 47.600 19.320 ;
      LAYER met1 ;
        RECT 47.600 18.760 47.880 19.320 ;
      LAYER met1 ;
        RECT 47.880 18.760 50.960 19.320 ;
      LAYER met1 ;
        RECT 50.960 19.040 51.240 19.320 ;
      LAYER met1 ;
        RECT 51.240 19.040 52.920 19.320 ;
      LAYER met1 ;
        RECT 52.920 19.040 54.320 19.320 ;
      LAYER met1 ;
        RECT 54.320 19.040 54.600 19.320 ;
      LAYER met1 ;
        RECT 54.600 19.040 54.880 19.600 ;
      LAYER met1 ;
        RECT 10.360 15.120 12.600 15.400 ;
      LAYER met1 ;
        RECT 12.600 15.120 14.000 15.400 ;
      LAYER met1 ;
        RECT 14.000 15.120 19.040 15.400 ;
        RECT 10.360 14.840 12.320 15.120 ;
      LAYER met1 ;
        RECT 12.320 14.840 13.720 15.120 ;
      LAYER met1 ;
        RECT 13.720 14.840 19.040 15.120 ;
      LAYER met1 ;
        RECT 19.040 14.840 20.440 15.400 ;
      LAYER met1 ;
        RECT 20.440 14.840 23.240 15.400 ;
      LAYER met1 ;
        RECT 23.240 15.120 26.600 15.400 ;
      LAYER met1 ;
        RECT 26.600 15.120 29.960 15.400 ;
      LAYER met1 ;
        RECT 23.240 14.840 26.040 15.120 ;
      LAYER met1 ;
        RECT 26.040 14.840 29.960 15.120 ;
      LAYER met1 ;
        RECT 29.960 14.840 31.360 15.400 ;
      LAYER met1 ;
        RECT 31.360 15.120 41.440 15.400 ;
      LAYER met1 ;
        RECT 41.440 15.120 43.120 15.400 ;
      LAYER met1 ;
        RECT 43.120 15.120 44.240 15.400 ;
      LAYER met1 ;
        RECT 44.240 15.120 44.520 15.400 ;
      LAYER met1 ;
        RECT 44.520 15.120 50.960 18.760 ;
      LAYER met1 ;
        RECT 50.960 15.120 51.520 19.040 ;
      LAYER met1 ;
        RECT 51.520 18.480 52.920 19.040 ;
      LAYER met1 ;
        RECT 52.920 18.760 54.880 19.040 ;
        RECT 52.920 18.480 53.760 18.760 ;
      LAYER met1 ;
        RECT 53.760 18.480 54.040 18.760 ;
      LAYER met1 ;
        RECT 54.040 18.480 54.880 18.760 ;
      LAYER met1 ;
        RECT 51.520 17.080 53.200 18.480 ;
      LAYER met1 ;
        RECT 53.200 17.080 53.760 18.480 ;
      LAYER met1 ;
        RECT 53.760 17.920 54.320 18.480 ;
      LAYER met1 ;
        RECT 54.320 17.920 54.880 18.480 ;
      LAYER met1 ;
        RECT 54.880 17.920 56.560 19.880 ;
      LAYER met1 ;
        RECT 56.560 18.200 57.120 20.160 ;
      LAYER met1 ;
        RECT 57.120 19.600 67.760 20.160 ;
      LAYER met1 ;
        RECT 67.760 19.880 72.240 20.720 ;
        RECT 67.760 19.600 69.720 19.880 ;
      LAYER met1 ;
        RECT 69.720 19.600 70.560 19.880 ;
        RECT 57.120 19.040 70.560 19.600 ;
      LAYER met1 ;
        RECT 70.560 19.320 72.240 19.880 ;
      LAYER met1 ;
        RECT 72.240 19.320 77.560 20.720 ;
      LAYER met1 ;
        RECT 70.560 19.040 74.200 19.320 ;
      LAYER met1 ;
        RECT 57.120 18.200 67.200 19.040 ;
      LAYER met1 ;
        RECT 56.560 17.920 57.400 18.200 ;
      LAYER met1 ;
        RECT 53.760 17.360 56.840 17.920 ;
      LAYER met1 ;
        RECT 56.840 17.360 57.400 17.920 ;
      LAYER met1 ;
        RECT 57.400 17.640 67.200 18.200 ;
      LAYER met1 ;
        RECT 67.200 17.640 74.200 19.040 ;
      LAYER met1 ;
        RECT 74.200 18.760 77.560 19.320 ;
      LAYER met1 ;
        RECT 77.560 18.760 79.240 21.280 ;
      LAYER met1 ;
        RECT 74.200 17.920 77.280 18.760 ;
      LAYER met1 ;
        RECT 77.280 18.200 79.240 18.760 ;
      LAYER met1 ;
        RECT 79.240 18.200 79.520 21.280 ;
      LAYER met1 ;
        RECT 77.280 17.920 78.960 18.200 ;
      LAYER met1 ;
        RECT 74.200 17.640 77.000 17.920 ;
        RECT 57.400 17.360 70.280 17.640 ;
        RECT 53.760 17.080 57.120 17.360 ;
        RECT 51.520 15.960 52.920 17.080 ;
      LAYER met1 ;
        RECT 52.920 15.960 53.480 17.080 ;
      LAYER met1 ;
        RECT 53.480 16.800 57.120 17.080 ;
      LAYER met1 ;
        RECT 57.120 16.800 57.680 17.360 ;
      LAYER met1 ;
        RECT 57.680 16.800 70.280 17.360 ;
      LAYER met1 ;
        RECT 70.280 17.080 72.240 17.640 ;
      LAYER met1 ;
        RECT 72.240 17.360 77.000 17.640 ;
      LAYER met1 ;
        RECT 77.000 17.360 78.960 17.920 ;
      LAYER met1 ;
        RECT 72.240 17.080 76.720 17.360 ;
      LAYER met1 ;
        RECT 76.720 17.080 78.960 17.360 ;
      LAYER met1 ;
        RECT 78.960 17.080 79.520 18.200 ;
      LAYER met1 ;
        RECT 79.520 17.080 81.200 21.560 ;
      LAYER met1 ;
        RECT 81.200 19.880 89.880 21.560 ;
      LAYER met1 ;
        RECT 89.880 19.880 91.840 21.560 ;
      LAYER met1 ;
        RECT 91.840 19.880 92.400 21.840 ;
        RECT 81.200 19.040 89.600 19.880 ;
      LAYER met1 ;
        RECT 89.600 19.040 91.560 19.880 ;
      LAYER met1 ;
        RECT 91.560 19.040 92.400 19.880 ;
        RECT 81.200 18.760 89.320 19.040 ;
        RECT 81.200 18.480 82.880 18.760 ;
      LAYER met1 ;
        RECT 82.880 18.480 83.440 18.760 ;
      LAYER met1 ;
        RECT 83.440 18.480 89.320 18.760 ;
      LAYER met1 ;
        RECT 89.320 18.480 91.280 19.040 ;
      LAYER met1 ;
        RECT 81.200 17.920 82.600 18.480 ;
      LAYER met1 ;
        RECT 82.600 18.200 83.720 18.480 ;
      LAYER met1 ;
        RECT 83.720 18.200 89.040 18.480 ;
      LAYER met1 ;
        RECT 89.040 18.200 91.280 18.480 ;
      LAYER met1 ;
        RECT 91.280 18.200 92.400 19.040 ;
      LAYER met1 ;
        RECT 82.600 17.920 84.280 18.200 ;
      LAYER met1 ;
        RECT 84.280 17.920 88.760 18.200 ;
      LAYER met1 ;
        RECT 88.760 17.920 91.000 18.200 ;
      LAYER met1 ;
        RECT 81.200 17.640 82.320 17.920 ;
      LAYER met1 ;
        RECT 82.320 17.640 84.560 17.920 ;
      LAYER met1 ;
        RECT 84.560 17.640 88.480 17.920 ;
      LAYER met1 ;
        RECT 88.480 17.640 91.000 17.920 ;
      LAYER met1 ;
        RECT 91.000 17.640 92.400 18.200 ;
        RECT 81.200 17.360 82.040 17.640 ;
      LAYER met1 ;
        RECT 82.040 17.360 84.560 17.640 ;
      LAYER met1 ;
        RECT 84.560 17.360 88.200 17.640 ;
      LAYER met1 ;
        RECT 88.200 17.360 90.720 17.640 ;
      LAYER met1 ;
        RECT 90.720 17.360 92.400 17.640 ;
        RECT 81.200 17.080 81.760 17.360 ;
      LAYER met1 ;
        RECT 81.760 17.080 84.280 17.360 ;
      LAYER met1 ;
        RECT 84.280 17.080 87.920 17.360 ;
      LAYER met1 ;
        RECT 87.920 17.080 90.440 17.360 ;
        RECT 70.280 16.800 71.960 17.080 ;
      LAYER met1 ;
        RECT 53.480 16.240 57.400 16.800 ;
      LAYER met1 ;
        RECT 57.400 16.240 57.960 16.800 ;
      LAYER met1 ;
        RECT 57.960 16.520 70.000 16.800 ;
      LAYER met1 ;
        RECT 70.000 16.520 71.960 16.800 ;
      LAYER met1 ;
        RECT 71.960 16.520 76.440 17.080 ;
      LAYER met1 ;
        RECT 76.440 16.800 78.680 17.080 ;
      LAYER met1 ;
        RECT 78.680 16.800 79.520 17.080 ;
      LAYER met1 ;
        RECT 79.520 16.800 84.000 17.080 ;
      LAYER met1 ;
        RECT 84.000 16.800 87.640 17.080 ;
      LAYER met1 ;
        RECT 87.640 16.800 90.440 17.080 ;
      LAYER met1 ;
        RECT 90.440 16.800 92.400 17.360 ;
      LAYER met1 ;
        RECT 76.440 16.520 78.400 16.800 ;
      LAYER met1 ;
        RECT 57.960 16.240 69.720 16.520 ;
      LAYER met1 ;
        RECT 69.720 16.240 71.680 16.520 ;
      LAYER met1 ;
        RECT 71.680 16.240 76.160 16.520 ;
      LAYER met1 ;
        RECT 76.160 16.240 78.400 16.520 ;
      LAYER met1 ;
        RECT 78.400 16.240 79.520 16.800 ;
      LAYER met1 ;
        RECT 79.520 16.520 83.720 16.800 ;
      LAYER met1 ;
        RECT 83.720 16.520 87.360 16.800 ;
      LAYER met1 ;
        RECT 87.360 16.520 90.160 16.800 ;
      LAYER met1 ;
        RECT 90.160 16.520 92.400 16.800 ;
      LAYER met1 ;
        RECT 79.520 16.240 83.440 16.520 ;
      LAYER met1 ;
        RECT 83.440 16.240 86.800 16.520 ;
      LAYER met1 ;
        RECT 86.800 16.240 89.880 16.520 ;
      LAYER met1 ;
        RECT 89.880 16.240 92.400 16.520 ;
        RECT 53.480 15.960 57.680 16.240 ;
        RECT 51.520 15.120 52.640 15.960 ;
        RECT 31.360 14.840 41.160 15.120 ;
      LAYER met1 ;
        RECT 41.160 14.840 42.000 15.120 ;
      LAYER met1 ;
        RECT 42.000 14.840 42.560 15.120 ;
      LAYER met1 ;
        RECT 42.560 14.840 43.400 15.120 ;
      LAYER met1 ;
        RECT 43.400 14.840 52.640 15.120 ;
        RECT 10.360 14.560 12.040 14.840 ;
      LAYER met1 ;
        RECT 12.040 14.560 13.720 14.840 ;
      LAYER met1 ;
        RECT 13.720 14.560 19.320 14.840 ;
      LAYER met1 ;
        RECT 19.320 14.560 20.720 14.840 ;
      LAYER met1 ;
        RECT 20.720 14.560 23.240 14.840 ;
      LAYER met1 ;
        RECT 23.240 14.560 25.480 14.840 ;
      LAYER met1 ;
        RECT 25.480 14.560 29.680 14.840 ;
      LAYER met1 ;
        RECT 29.680 14.560 31.080 14.840 ;
      LAYER met1 ;
        RECT 31.080 14.560 41.160 14.840 ;
      LAYER met1 ;
        RECT 41.160 14.560 41.720 14.840 ;
      LAYER met1 ;
        RECT 10.360 14.280 11.760 14.560 ;
      LAYER met1 ;
        RECT 11.760 14.280 13.440 14.560 ;
      LAYER met1 ;
        RECT 13.440 14.280 19.600 14.560 ;
      LAYER met1 ;
        RECT 19.600 14.280 21.000 14.560 ;
      LAYER met1 ;
        RECT 21.000 14.280 29.400 14.560 ;
      LAYER met1 ;
        RECT 29.400 14.280 31.080 14.560 ;
      LAYER met1 ;
        RECT 31.080 14.280 40.880 14.560 ;
      LAYER met1 ;
        RECT 40.880 14.280 41.720 14.560 ;
      LAYER met1 ;
        RECT 41.720 14.280 42.560 14.840 ;
      LAYER met1 ;
        RECT 42.560 14.560 43.680 14.840 ;
      LAYER met1 ;
        RECT 43.680 14.560 52.640 14.840 ;
      LAYER met1 ;
        RECT 52.640 14.560 53.200 15.960 ;
      LAYER met1 ;
        RECT 53.200 15.680 57.680 15.960 ;
        RECT 53.200 14.560 55.440 15.680 ;
      LAYER met1 ;
        RECT 55.440 15.120 55.720 15.680 ;
      LAYER met1 ;
        RECT 55.720 15.400 57.680 15.680 ;
        RECT 55.720 15.120 56.840 15.400 ;
      LAYER met1 ;
        RECT 56.840 15.120 57.120 15.400 ;
      LAYER met1 ;
        RECT 57.120 15.120 57.680 15.400 ;
      LAYER met1 ;
        RECT 42.560 14.280 43.960 14.560 ;
      LAYER met1 ;
        RECT 43.960 14.280 46.200 14.560 ;
        RECT 10.360 14.000 11.480 14.280 ;
      LAYER met1 ;
        RECT 11.480 14.000 13.160 14.280 ;
      LAYER met1 ;
        RECT 13.160 14.000 19.600 14.280 ;
      LAYER met1 ;
        RECT 19.600 14.000 21.280 14.280 ;
      LAYER met1 ;
        RECT 21.280 14.000 29.120 14.280 ;
      LAYER met1 ;
        RECT 29.120 14.000 30.800 14.280 ;
      LAYER met1 ;
        RECT 30.800 14.000 40.880 14.280 ;
        RECT 10.360 13.720 11.200 14.000 ;
      LAYER met1 ;
        RECT 11.200 13.720 12.880 14.000 ;
      LAYER met1 ;
        RECT 12.880 13.720 19.880 14.000 ;
      LAYER met1 ;
        RECT 19.880 13.720 21.560 14.000 ;
      LAYER met1 ;
        RECT 21.560 13.720 28.840 14.000 ;
      LAYER met1 ;
        RECT 28.840 13.720 30.520 14.000 ;
      LAYER met1 ;
        RECT 30.520 13.720 40.880 14.000 ;
      LAYER met1 ;
        RECT 40.880 13.720 42.280 14.280 ;
      LAYER met1 ;
        RECT 42.280 13.720 42.560 14.280 ;
      LAYER met1 ;
        RECT 42.560 13.720 43.120 14.280 ;
      LAYER met1 ;
        RECT 43.120 14.000 43.400 14.280 ;
      LAYER met1 ;
        RECT 43.400 14.000 44.520 14.280 ;
      LAYER met1 ;
        RECT 44.520 14.000 46.200 14.280 ;
      LAYER met1 ;
        RECT 46.200 14.000 50.400 14.560 ;
      LAYER met1 ;
        RECT 50.400 14.280 52.640 14.560 ;
      LAYER met1 ;
        RECT 52.640 14.280 53.480 14.560 ;
      LAYER met1 ;
        RECT 43.120 13.720 43.680 14.000 ;
      LAYER met1 ;
        RECT 43.680 13.720 44.800 14.000 ;
      LAYER met1 ;
        RECT 44.800 13.720 46.200 14.000 ;
      LAYER met1 ;
        RECT 46.200 13.720 46.760 14.000 ;
      LAYER met1 ;
        RECT 46.760 13.720 49.840 14.000 ;
        RECT 0.000 12.320 4.200 12.600 ;
      LAYER met1 ;
        RECT 4.200 12.320 10.360 12.600 ;
      LAYER met1 ;
        RECT 10.360 12.320 10.920 13.720 ;
      LAYER met1 ;
        RECT 10.920 13.440 12.600 13.720 ;
      LAYER met1 ;
        RECT 12.600 13.440 20.160 13.720 ;
      LAYER met1 ;
        RECT 20.160 13.440 22.120 13.720 ;
      LAYER met1 ;
        RECT 22.120 13.440 28.280 13.720 ;
      LAYER met1 ;
        RECT 28.280 13.440 30.240 13.720 ;
      LAYER met1 ;
        RECT 30.240 13.440 41.160 13.720 ;
      LAYER met1 ;
        RECT 41.160 13.440 43.120 13.720 ;
      LAYER met1 ;
        RECT 43.120 13.440 43.400 13.720 ;
      LAYER met1 ;
        RECT 43.400 13.440 45.640 13.720 ;
      LAYER met1 ;
        RECT 45.640 13.440 46.480 13.720 ;
      LAYER met1 ;
        RECT 10.920 13.160 12.320 13.440 ;
      LAYER met1 ;
        RECT 12.320 13.160 20.440 13.440 ;
      LAYER met1 ;
        RECT 20.440 13.160 22.680 13.440 ;
      LAYER met1 ;
        RECT 22.680 13.160 27.720 13.440 ;
      LAYER met1 ;
        RECT 27.720 13.160 29.960 13.440 ;
      LAYER met1 ;
        RECT 29.960 13.160 41.440 13.440 ;
      LAYER met1 ;
        RECT 41.440 13.160 46.200 13.440 ;
      LAYER met1 ;
        RECT 46.200 13.160 46.480 13.440 ;
      LAYER met1 ;
        RECT 46.480 13.160 47.040 13.720 ;
      LAYER met1 ;
        RECT 47.040 13.160 49.840 13.720 ;
      LAYER met1 ;
        RECT 10.920 12.880 12.040 13.160 ;
      LAYER met1 ;
        RECT 12.040 12.880 20.720 13.160 ;
      LAYER met1 ;
        RECT 20.720 12.880 23.240 13.160 ;
      LAYER met1 ;
        RECT 23.240 12.880 27.160 13.160 ;
      LAYER met1 ;
        RECT 27.160 12.880 29.680 13.160 ;
      LAYER met1 ;
        RECT 29.680 12.880 41.440 13.160 ;
      LAYER met1 ;
        RECT 41.440 12.880 47.320 13.160 ;
      LAYER met1 ;
        RECT 47.320 12.880 49.840 13.160 ;
      LAYER met1 ;
        RECT 49.840 12.880 50.400 14.000 ;
      LAYER met1 ;
        RECT 50.400 13.720 52.920 14.280 ;
      LAYER met1 ;
        RECT 52.920 13.720 53.480 14.280 ;
      LAYER met1 ;
        RECT 50.400 13.440 52.640 13.720 ;
      LAYER met1 ;
        RECT 52.640 13.440 53.480 13.720 ;
      LAYER met1 ;
        RECT 50.400 13.160 52.360 13.440 ;
      LAYER met1 ;
        RECT 52.360 13.160 53.480 13.440 ;
      LAYER met1 ;
        RECT 53.480 13.160 53.760 14.560 ;
      LAYER met1 ;
        RECT 53.760 14.280 54.320 14.560 ;
      LAYER met1 ;
        RECT 54.320 14.280 55.440 14.560 ;
      LAYER met1 ;
        RECT 53.760 13.160 54.880 14.280 ;
      LAYER met1 ;
        RECT 54.880 13.440 55.440 14.280 ;
      LAYER met1 ;
        RECT 55.440 13.720 56.000 15.120 ;
      LAYER met1 ;
        RECT 56.000 14.560 56.840 15.120 ;
      LAYER met1 ;
        RECT 56.840 14.840 57.400 15.120 ;
      LAYER met1 ;
        RECT 57.400 14.840 57.680 15.120 ;
      LAYER met1 ;
        RECT 57.680 14.840 58.240 16.240 ;
      LAYER met1 ;
        RECT 58.240 15.960 69.440 16.240 ;
      LAYER met1 ;
        RECT 69.440 15.960 71.680 16.240 ;
      LAYER met1 ;
        RECT 71.680 15.960 75.880 16.240 ;
        RECT 58.240 15.120 68.880 15.960 ;
      LAYER met1 ;
        RECT 68.880 15.680 71.400 15.960 ;
      LAYER met1 ;
        RECT 71.400 15.680 75.880 15.960 ;
      LAYER met1 ;
        RECT 75.880 15.680 78.120 16.240 ;
      LAYER met1 ;
        RECT 78.120 15.680 79.520 16.240 ;
      LAYER met1 ;
        RECT 79.520 15.960 83.160 16.240 ;
      LAYER met1 ;
        RECT 83.160 15.960 86.240 16.240 ;
      LAYER met1 ;
        RECT 86.240 15.960 89.600 16.240 ;
      LAYER met1 ;
        RECT 89.600 15.960 92.400 16.240 ;
      LAYER met1 ;
        RECT 79.520 15.680 82.880 15.960 ;
      LAYER met1 ;
        RECT 82.880 15.680 85.680 15.960 ;
      LAYER met1 ;
        RECT 85.680 15.680 89.320 15.960 ;
      LAYER met1 ;
        RECT 89.320 15.680 92.400 15.960 ;
      LAYER met1 ;
        RECT 68.880 15.400 71.120 15.680 ;
      LAYER met1 ;
        RECT 71.120 15.400 76.160 15.680 ;
      LAYER met1 ;
        RECT 76.160 15.400 77.840 15.680 ;
      LAYER met1 ;
        RECT 77.840 15.400 79.520 15.680 ;
      LAYER met1 ;
        RECT 79.520 15.400 82.320 15.680 ;
      LAYER met1 ;
        RECT 82.320 15.400 85.680 15.680 ;
      LAYER met1 ;
        RECT 85.680 15.400 88.760 15.680 ;
      LAYER met1 ;
        RECT 88.760 15.400 92.400 15.680 ;
      LAYER met1 ;
        RECT 68.880 15.120 70.840 15.400 ;
      LAYER met1 ;
        RECT 70.840 15.120 76.440 15.400 ;
      LAYER met1 ;
        RECT 76.440 15.120 77.560 15.400 ;
      LAYER met1 ;
        RECT 77.560 15.120 79.520 15.400 ;
      LAYER met1 ;
        RECT 79.520 15.120 81.760 15.400 ;
      LAYER met1 ;
        RECT 81.760 15.120 85.960 15.400 ;
      LAYER met1 ;
        RECT 85.960 15.120 88.200 15.400 ;
      LAYER met1 ;
        RECT 88.200 15.120 92.400 15.400 ;
        RECT 58.240 14.840 69.160 15.120 ;
      LAYER met1 ;
        RECT 69.160 14.840 70.560 15.120 ;
      LAYER met1 ;
        RECT 70.560 14.840 76.440 15.120 ;
      LAYER met1 ;
        RECT 76.440 14.840 77.000 15.120 ;
      LAYER met1 ;
        RECT 77.000 14.840 80.080 15.120 ;
      LAYER met1 ;
        RECT 80.080 14.840 80.920 15.120 ;
      LAYER met1 ;
        RECT 80.920 14.840 86.240 15.120 ;
      LAYER met1 ;
        RECT 86.240 14.840 87.640 15.120 ;
      LAYER met1 ;
        RECT 87.640 14.840 92.400 15.120 ;
      LAYER met1 ;
        RECT 56.840 14.560 58.240 14.840 ;
      LAYER met1 ;
        RECT 58.240 14.560 69.440 14.840 ;
      LAYER met1 ;
        RECT 69.440 14.560 70.000 14.840 ;
      LAYER met1 ;
        RECT 70.000 14.560 92.400 14.840 ;
        RECT 56.000 14.000 57.120 14.560 ;
      LAYER met1 ;
        RECT 57.120 14.000 59.080 14.560 ;
      LAYER met1 ;
        RECT 59.080 14.000 92.400 14.560 ;
        RECT 56.000 13.720 56.280 14.000 ;
      LAYER met1 ;
        RECT 56.280 13.720 56.840 14.000 ;
      LAYER met1 ;
        RECT 56.840 13.720 57.120 14.000 ;
      LAYER met1 ;
        RECT 57.120 13.720 57.680 14.000 ;
      LAYER met1 ;
        RECT 57.680 13.720 58.240 14.000 ;
      LAYER met1 ;
        RECT 58.240 13.720 58.800 14.000 ;
      LAYER met1 ;
        RECT 58.800 13.720 92.400 14.000 ;
      LAYER met1 ;
        RECT 55.440 13.440 55.720 13.720 ;
      LAYER met1 ;
        RECT 54.880 13.160 55.160 13.440 ;
      LAYER met1 ;
        RECT 55.160 13.160 55.720 13.440 ;
      LAYER met1 ;
        RECT 50.400 12.880 52.080 13.160 ;
      LAYER met1 ;
        RECT 52.080 12.880 55.720 13.160 ;
      LAYER met1 ;
        RECT 55.720 12.880 56.280 13.720 ;
      LAYER met1 ;
        RECT 56.280 13.440 57.400 13.720 ;
      LAYER met1 ;
        RECT 57.400 13.440 57.960 13.720 ;
      LAYER met1 ;
        RECT 57.960 13.440 58.520 13.720 ;
      LAYER met1 ;
        RECT 58.520 13.440 92.400 13.720 ;
      LAYER met1 ;
        RECT 56.280 12.880 57.120 13.440 ;
      LAYER met1 ;
        RECT 57.120 13.160 57.680 13.440 ;
      LAYER met1 ;
        RECT 57.680 13.160 58.240 13.440 ;
      LAYER met1 ;
        RECT 58.240 13.160 92.400 13.440 ;
        RECT 57.120 12.880 57.400 13.160 ;
      LAYER met1 ;
        RECT 10.920 12.600 11.760 12.880 ;
      LAYER met1 ;
        RECT 11.760 12.600 21.280 12.880 ;
      LAYER met1 ;
        RECT 21.280 12.600 24.360 12.880 ;
      LAYER met1 ;
        RECT 24.360 12.600 26.040 12.880 ;
      LAYER met1 ;
        RECT 26.040 12.600 29.120 12.880 ;
      LAYER met1 ;
        RECT 29.120 12.600 41.720 12.880 ;
      LAYER met1 ;
        RECT 41.720 12.600 45.640 12.880 ;
      LAYER met1 ;
        RECT 45.640 12.600 45.920 12.880 ;
      LAYER met1 ;
        RECT 45.920 12.600 47.600 12.880 ;
      LAYER met1 ;
        RECT 47.600 12.600 49.560 12.880 ;
      LAYER met1 ;
        RECT 49.560 12.600 50.120 12.880 ;
      LAYER met1 ;
        RECT 50.120 12.600 51.240 12.880 ;
      LAYER met1 ;
        RECT 51.240 12.600 55.720 12.880 ;
      LAYER met1 ;
        RECT 55.720 12.600 56.000 12.880 ;
      LAYER met1 ;
        RECT 56.000 12.600 56.840 12.880 ;
      LAYER met1 ;
        RECT 56.840 12.600 57.400 12.880 ;
      LAYER met1 ;
        RECT 57.400 12.600 57.960 13.160 ;
      LAYER met1 ;
        RECT 57.960 12.600 92.400 13.160 ;
      LAYER met1 ;
        RECT 10.920 12.320 11.480 12.600 ;
      LAYER met1 ;
        RECT 11.480 12.320 21.560 12.600 ;
      LAYER met1 ;
        RECT 21.560 12.320 28.840 12.600 ;
      LAYER met1 ;
        RECT 28.840 12.320 42.280 12.600 ;
      LAYER met1 ;
        RECT 42.280 12.320 42.840 12.600 ;
      LAYER met1 ;
        RECT 42.840 12.320 43.400 12.600 ;
      LAYER met1 ;
        RECT 43.400 12.320 43.960 12.600 ;
      LAYER met1 ;
        RECT 43.960 12.320 44.800 12.600 ;
      LAYER met1 ;
        RECT 44.800 12.320 45.360 12.600 ;
      LAYER met1 ;
        RECT 45.360 12.320 46.200 12.600 ;
      LAYER met1 ;
        RECT 46.200 12.320 52.360 12.600 ;
      LAYER met1 ;
        RECT 52.360 12.320 52.640 12.600 ;
      LAYER met1 ;
        RECT 52.640 12.320 56.560 12.600 ;
      LAYER met1 ;
        RECT 56.560 12.320 57.120 12.600 ;
      LAYER met1 ;
        RECT 57.120 12.320 57.680 12.600 ;
      LAYER met1 ;
        RECT 57.680 12.320 92.400 12.600 ;
        RECT 0.000 12.040 4.760 12.320 ;
      LAYER met1 ;
        RECT 4.760 12.040 10.360 12.320 ;
      LAYER met1 ;
        RECT 10.360 12.040 22.120 12.320 ;
      LAYER met1 ;
        RECT 22.120 12.040 28.280 12.320 ;
      LAYER met1 ;
        RECT 28.280 12.040 42.560 12.320 ;
      LAYER met1 ;
        RECT 42.560 12.040 43.120 12.320 ;
      LAYER met1 ;
        RECT 43.120 12.040 46.200 12.320 ;
      LAYER met1 ;
        RECT 46.200 12.040 47.040 12.320 ;
      LAYER met1 ;
        RECT 47.040 12.040 47.600 12.320 ;
        RECT 0.000 11.760 5.320 12.040 ;
      LAYER met1 ;
        RECT 5.320 11.760 10.080 12.040 ;
      LAYER met1 ;
        RECT 10.080 11.760 22.680 12.040 ;
      LAYER met1 ;
        RECT 22.680 11.760 27.720 12.040 ;
      LAYER met1 ;
        RECT 27.720 11.760 42.560 12.040 ;
      LAYER met1 ;
        RECT 42.560 11.760 43.400 12.040 ;
      LAYER met1 ;
        RECT 43.400 11.760 46.480 12.040 ;
      LAYER met1 ;
        RECT 46.480 11.760 47.320 12.040 ;
      LAYER met1 ;
        RECT 47.320 11.760 47.600 12.040 ;
      LAYER met1 ;
        RECT 47.600 11.760 52.080 12.320 ;
      LAYER met1 ;
        RECT 52.080 12.040 52.920 12.320 ;
      LAYER met1 ;
        RECT 52.920 12.040 53.480 12.320 ;
      LAYER met1 ;
        RECT 53.480 12.040 54.040 12.320 ;
      LAYER met1 ;
        RECT 54.040 12.040 54.880 12.320 ;
      LAYER met1 ;
        RECT 54.880 12.040 55.160 12.320 ;
      LAYER met1 ;
        RECT 55.160 12.040 55.720 12.320 ;
      LAYER met1 ;
        RECT 55.720 12.040 56.840 12.320 ;
      LAYER met1 ;
        RECT 56.840 12.040 57.400 12.320 ;
      LAYER met1 ;
        RECT 57.400 12.040 92.400 12.320 ;
        RECT 52.080 11.760 52.640 12.040 ;
      LAYER met1 ;
        RECT 52.640 11.760 53.480 12.040 ;
      LAYER met1 ;
        RECT 53.480 11.760 56.560 12.040 ;
      LAYER met1 ;
        RECT 56.560 11.760 57.120 12.040 ;
      LAYER met1 ;
        RECT 57.120 11.760 92.400 12.040 ;
        RECT 0.000 11.480 6.160 11.760 ;
      LAYER met1 ;
        RECT 6.160 11.480 9.240 11.760 ;
      LAYER met1 ;
        RECT 9.240 11.480 23.800 11.760 ;
      LAYER met1 ;
        RECT 23.800 11.480 26.600 11.760 ;
      LAYER met1 ;
        RECT 26.600 11.480 42.840 11.760 ;
      LAYER met1 ;
        RECT 42.840 11.480 43.680 11.760 ;
      LAYER met1 ;
        RECT 43.680 11.480 46.760 11.760 ;
      LAYER met1 ;
        RECT 46.760 11.480 49.280 11.760 ;
      LAYER met1 ;
        RECT 0.000 11.200 43.120 11.480 ;
      LAYER met1 ;
        RECT 43.120 11.200 43.960 11.480 ;
      LAYER met1 ;
        RECT 43.960 11.200 47.040 11.480 ;
      LAYER met1 ;
        RECT 47.040 11.200 49.280 11.480 ;
      LAYER met1 ;
        RECT 49.280 11.200 49.560 11.760 ;
      LAYER met1 ;
        RECT 49.560 11.480 50.120 11.760 ;
      LAYER met1 ;
        RECT 50.120 11.480 50.680 11.760 ;
      LAYER met1 ;
        RECT 50.680 11.480 52.920 11.760 ;
      LAYER met1 ;
        RECT 52.920 11.480 53.200 11.760 ;
      LAYER met1 ;
        RECT 53.200 11.480 53.480 11.760 ;
      LAYER met1 ;
        RECT 53.480 11.480 56.280 11.760 ;
      LAYER met1 ;
        RECT 56.280 11.480 56.840 11.760 ;
      LAYER met1 ;
        RECT 56.840 11.480 92.400 11.760 ;
      LAYER met1 ;
        RECT 49.560 11.200 50.960 11.480 ;
      LAYER met1 ;
        RECT 0.000 10.920 43.400 11.200 ;
      LAYER met1 ;
        RECT 43.400 10.920 45.080 11.200 ;
      LAYER met1 ;
        RECT 45.080 10.920 47.040 11.200 ;
        RECT 0.000 10.640 43.680 10.920 ;
      LAYER met1 ;
        RECT 43.680 10.640 46.760 10.920 ;
      LAYER met1 ;
        RECT 46.760 10.640 47.040 10.920 ;
      LAYER met1 ;
        RECT 47.040 10.640 50.400 11.200 ;
      LAYER met1 ;
        RECT 50.400 10.640 50.680 11.200 ;
      LAYER met1 ;
        RECT 50.680 10.640 50.960 11.200 ;
      LAYER met1 ;
        RECT 0.000 10.360 45.080 10.640 ;
      LAYER met1 ;
        RECT 45.080 10.360 47.600 10.640 ;
      LAYER met1 ;
        RECT 47.600 10.360 47.880 10.640 ;
        RECT 0.000 9.800 46.480 10.360 ;
      LAYER met1 ;
        RECT 46.480 9.800 47.320 10.360 ;
      LAYER met1 ;
        RECT 47.320 10.080 47.880 10.360 ;
      LAYER met1 ;
        RECT 47.880 10.080 48.440 10.640 ;
      LAYER met1 ;
        RECT 48.440 10.080 49.000 10.640 ;
      LAYER met1 ;
        RECT 49.000 10.360 50.960 10.640 ;
      LAYER met1 ;
        RECT 50.960 10.360 51.240 11.480 ;
      LAYER met1 ;
        RECT 51.240 10.920 52.640 11.480 ;
      LAYER met1 ;
        RECT 52.640 11.200 56.000 11.480 ;
      LAYER met1 ;
        RECT 56.000 11.200 56.560 11.480 ;
      LAYER met1 ;
        RECT 56.560 11.200 92.400 11.480 ;
        RECT 52.640 10.920 54.880 11.200 ;
      LAYER met1 ;
        RECT 54.880 10.920 56.280 11.200 ;
      LAYER met1 ;
        RECT 56.280 10.920 92.400 11.200 ;
      LAYER met1 ;
        RECT 51.240 10.640 52.920 10.920 ;
      LAYER met1 ;
        RECT 52.920 10.640 53.200 10.920 ;
      LAYER met1 ;
        RECT 53.200 10.640 56.000 10.920 ;
      LAYER met1 ;
        RECT 56.000 10.640 92.400 10.920 ;
      LAYER met1 ;
        RECT 51.240 10.360 52.080 10.640 ;
        RECT 49.000 10.080 50.680 10.360 ;
      LAYER met1 ;
        RECT 50.680 10.080 51.520 10.360 ;
      LAYER met1 ;
        RECT 51.520 10.080 52.080 10.360 ;
      LAYER met1 ;
        RECT 52.080 10.080 52.360 10.640 ;
      LAYER met1 ;
        RECT 52.360 10.360 54.880 10.640 ;
      LAYER met1 ;
        RECT 54.880 10.360 92.400 10.640 ;
      LAYER met1 ;
        RECT 52.360 10.080 53.200 10.360 ;
      LAYER met1 ;
        RECT 47.320 9.800 47.600 10.080 ;
      LAYER met1 ;
        RECT 47.600 9.800 48.440 10.080 ;
      LAYER met1 ;
        RECT 48.440 9.800 49.560 10.080 ;
      LAYER met1 ;
        RECT 49.560 9.800 50.120 10.080 ;
      LAYER met1 ;
        RECT 50.120 9.800 51.520 10.080 ;
      LAYER met1 ;
        RECT 51.520 9.800 53.200 10.080 ;
      LAYER met1 ;
        RECT 53.200 9.800 92.400 10.360 ;
        RECT 0.000 9.520 46.760 9.800 ;
        RECT 0.000 9.240 43.400 9.520 ;
      LAYER met1 ;
        RECT 43.400 9.240 44.240 9.520 ;
      LAYER met1 ;
        RECT 44.240 9.240 46.760 9.520 ;
      LAYER met1 ;
        RECT 46.760 9.240 48.160 9.800 ;
      LAYER met1 ;
        RECT 0.000 8.960 42.560 9.240 ;
      LAYER met1 ;
        RECT 42.560 8.960 44.800 9.240 ;
      LAYER met1 ;
        RECT 44.800 8.960 46.480 9.240 ;
      LAYER met1 ;
        RECT 46.480 8.960 48.160 9.240 ;
      LAYER met1 ;
        RECT 48.160 8.960 51.520 9.800 ;
      LAYER met1 ;
        RECT 51.520 9.520 52.920 9.800 ;
      LAYER met1 ;
        RECT 52.920 9.520 92.400 9.800 ;
      LAYER met1 ;
        RECT 51.520 8.960 53.200 9.520 ;
      LAYER met1 ;
        RECT 53.200 9.240 54.880 9.520 ;
      LAYER met1 ;
        RECT 54.880 9.240 56.000 9.520 ;
      LAYER met1 ;
        RECT 56.000 9.240 92.400 9.520 ;
        RECT 53.200 8.960 54.320 9.240 ;
      LAYER met1 ;
        RECT 54.320 8.960 57.120 9.240 ;
      LAYER met1 ;
        RECT 57.120 8.960 92.400 9.240 ;
        RECT 0.000 8.680 41.440 8.960 ;
      LAYER met1 ;
        RECT 41.440 8.680 43.400 8.960 ;
      LAYER met1 ;
        RECT 43.400 8.680 44.240 8.960 ;
      LAYER met1 ;
        RECT 44.240 8.680 45.360 8.960 ;
      LAYER met1 ;
        RECT 45.360 8.680 46.480 8.960 ;
      LAYER met1 ;
        RECT 46.480 8.680 47.880 8.960 ;
      LAYER met1 ;
        RECT 0.000 8.400 40.320 8.680 ;
      LAYER met1 ;
        RECT 40.320 8.400 42.560 8.680 ;
      LAYER met1 ;
        RECT 42.560 8.400 44.800 8.680 ;
      LAYER met1 ;
        RECT 44.800 8.400 45.920 8.680 ;
      LAYER met1 ;
        RECT 45.920 8.400 46.200 8.680 ;
      LAYER met1 ;
        RECT 46.200 8.400 47.040 8.680 ;
      LAYER met1 ;
        RECT 47.040 8.400 47.320 8.680 ;
        RECT 0.000 7.840 39.760 8.400 ;
      LAYER met1 ;
        RECT 39.760 8.120 41.440 8.400 ;
      LAYER met1 ;
        RECT 41.440 8.120 45.360 8.400 ;
      LAYER met1 ;
        RECT 45.360 8.120 46.760 8.400 ;
      LAYER met1 ;
        RECT 46.760 8.120 47.320 8.400 ;
      LAYER met1 ;
        RECT 47.320 8.120 47.880 8.680 ;
      LAYER met1 ;
        RECT 47.880 8.120 51.800 8.960 ;
      LAYER met1 ;
        RECT 51.800 8.680 53.200 8.960 ;
      LAYER met1 ;
        RECT 53.200 8.680 53.760 8.960 ;
      LAYER met1 ;
        RECT 53.760 8.680 54.880 8.960 ;
      LAYER met1 ;
        RECT 54.880 8.680 56.000 8.960 ;
      LAYER met1 ;
        RECT 56.000 8.680 57.960 8.960 ;
      LAYER met1 ;
        RECT 57.960 8.680 92.400 8.960 ;
      LAYER met1 ;
        RECT 39.760 7.840 40.600 8.120 ;
      LAYER met1 ;
        RECT 40.600 7.840 45.920 8.120 ;
        RECT 0.000 7.560 40.040 7.840 ;
      LAYER met1 ;
        RECT 40.040 7.560 41.160 7.840 ;
      LAYER met1 ;
        RECT 41.160 7.560 45.920 7.840 ;
      LAYER met1 ;
        RECT 45.920 7.560 46.760 8.120 ;
      LAYER met1 ;
        RECT 46.760 7.560 47.040 8.120 ;
        RECT 0.000 7.280 40.600 7.560 ;
      LAYER met1 ;
        RECT 40.600 7.280 41.720 7.560 ;
      LAYER met1 ;
        RECT 41.720 7.280 45.920 7.560 ;
      LAYER met1 ;
        RECT 45.920 7.280 46.480 7.560 ;
      LAYER met1 ;
        RECT 46.480 7.280 47.040 7.560 ;
      LAYER met1 ;
        RECT 47.040 7.280 47.600 8.120 ;
      LAYER met1 ;
        RECT 47.600 7.560 51.800 8.120 ;
      LAYER met1 ;
        RECT 51.800 7.840 52.360 8.680 ;
      LAYER met1 ;
        RECT 52.360 8.120 52.640 8.680 ;
      LAYER met1 ;
        RECT 52.640 8.400 54.320 8.680 ;
      LAYER met1 ;
        RECT 54.320 8.400 57.120 8.680 ;
      LAYER met1 ;
        RECT 57.120 8.400 59.080 8.680 ;
      LAYER met1 ;
        RECT 59.080 8.400 92.400 8.680 ;
      LAYER met1 ;
        RECT 52.640 8.120 54.040 8.400 ;
      LAYER met1 ;
        RECT 54.040 8.120 57.960 8.400 ;
      LAYER met1 ;
        RECT 57.960 8.120 59.640 8.400 ;
      LAYER met1 ;
        RECT 52.360 7.840 52.920 8.120 ;
      LAYER met1 ;
        RECT 52.920 7.840 53.480 8.120 ;
      LAYER met1 ;
        RECT 53.480 7.840 58.800 8.120 ;
      LAYER met1 ;
        RECT 58.800 7.840 59.640 8.120 ;
      LAYER met1 ;
        RECT 59.640 7.840 92.400 8.400 ;
      LAYER met1 ;
        RECT 51.800 7.560 52.640 7.840 ;
      LAYER met1 ;
        RECT 47.600 7.280 52.080 7.560 ;
        RECT 0.000 7.000 41.160 7.280 ;
      LAYER met1 ;
        RECT 41.160 7.000 42.280 7.280 ;
      LAYER met1 ;
        RECT 42.280 7.000 45.640 7.280 ;
      LAYER met1 ;
        RECT 45.640 7.000 46.480 7.280 ;
      LAYER met1 ;
        RECT 46.480 7.000 46.760 7.280 ;
        RECT 0.000 6.720 41.720 7.000 ;
      LAYER met1 ;
        RECT 41.720 6.720 42.840 7.000 ;
      LAYER met1 ;
        RECT 42.840 6.720 45.640 7.000 ;
      LAYER met1 ;
        RECT 45.640 6.720 46.200 7.000 ;
      LAYER met1 ;
        RECT 46.200 6.720 46.760 7.000 ;
      LAYER met1 ;
        RECT 46.760 6.720 47.320 7.280 ;
      LAYER met1 ;
        RECT 0.000 6.440 42.280 6.720 ;
      LAYER met1 ;
        RECT 42.280 6.440 43.400 6.720 ;
      LAYER met1 ;
        RECT 43.400 6.440 44.520 6.720 ;
      LAYER met1 ;
        RECT 44.520 6.440 46.200 6.720 ;
      LAYER met1 ;
        RECT 46.200 6.440 46.480 6.720 ;
      LAYER met1 ;
        RECT 46.480 6.440 47.320 6.720 ;
      LAYER met1 ;
        RECT 47.320 6.440 52.080 7.280 ;
      LAYER met1 ;
        RECT 52.080 7.000 52.640 7.560 ;
      LAYER met1 ;
        RECT 52.640 7.280 52.920 7.840 ;
      LAYER met1 ;
        RECT 52.920 7.280 53.760 7.840 ;
      LAYER met1 ;
        RECT 53.760 7.560 58.240 7.840 ;
      LAYER met1 ;
        RECT 58.240 7.560 59.360 7.840 ;
      LAYER met1 ;
        RECT 59.360 7.560 92.400 7.840 ;
        RECT 53.760 7.280 57.680 7.560 ;
      LAYER met1 ;
        RECT 57.680 7.280 58.800 7.560 ;
      LAYER met1 ;
        RECT 58.800 7.280 92.400 7.560 ;
        RECT 52.640 7.000 53.200 7.280 ;
      LAYER met1 ;
        RECT 53.200 7.000 53.760 7.280 ;
      LAYER met1 ;
        RECT 53.760 7.000 57.120 7.280 ;
      LAYER met1 ;
        RECT 57.120 7.000 58.240 7.280 ;
      LAYER met1 ;
        RECT 58.240 7.000 92.400 7.280 ;
        RECT 0.000 6.160 42.840 6.440 ;
      LAYER met1 ;
        RECT 42.840 6.160 47.040 6.440 ;
      LAYER met1 ;
        RECT 0.000 5.880 43.400 6.160 ;
      LAYER met1 ;
        RECT 43.400 5.880 44.520 6.160 ;
      LAYER met1 ;
        RECT 44.520 5.880 45.640 6.160 ;
      LAYER met1 ;
        RECT 45.640 5.880 47.040 6.160 ;
      LAYER met1 ;
        RECT 47.040 5.880 52.080 6.440 ;
      LAYER met1 ;
        RECT 52.080 6.160 52.920 7.000 ;
      LAYER met1 ;
        RECT 52.920 6.160 53.200 7.000 ;
      LAYER met1 ;
        RECT 53.200 6.720 54.040 7.000 ;
      LAYER met1 ;
        RECT 54.040 6.720 56.560 7.000 ;
      LAYER met1 ;
        RECT 56.560 6.720 57.680 7.000 ;
      LAYER met1 ;
        RECT 57.680 6.720 92.400 7.000 ;
      LAYER met1 ;
        RECT 53.200 6.440 54.880 6.720 ;
      LAYER met1 ;
        RECT 54.880 6.440 56.000 6.720 ;
      LAYER met1 ;
        RECT 56.000 6.440 57.120 6.720 ;
      LAYER met1 ;
        RECT 57.120 6.440 92.400 6.720 ;
      LAYER met1 ;
        RECT 53.200 6.160 56.560 6.440 ;
      LAYER met1 ;
        RECT 56.560 6.160 92.400 6.440 ;
      LAYER met1 ;
        RECT 52.080 5.880 54.040 6.160 ;
      LAYER met1 ;
        RECT 54.040 5.880 54.880 6.160 ;
      LAYER met1 ;
        RECT 54.880 5.880 56.000 6.160 ;
      LAYER met1 ;
        RECT 56.000 5.880 92.400 6.160 ;
        RECT 0.000 5.040 46.200 5.880 ;
      LAYER met1 ;
        RECT 46.200 5.600 47.040 5.880 ;
      LAYER met1 ;
        RECT 47.040 5.600 52.360 5.880 ;
      LAYER met1 ;
        RECT 52.360 5.600 54.040 5.880 ;
      LAYER met1 ;
        RECT 54.040 5.600 92.400 5.880 ;
      LAYER met1 ;
        RECT 46.200 5.040 46.760 5.600 ;
      LAYER met1 ;
        RECT 46.760 5.040 52.360 5.600 ;
        RECT 0.000 4.760 45.920 5.040 ;
      LAYER met1 ;
        RECT 45.920 4.760 46.480 5.040 ;
      LAYER met1 ;
        RECT 0.000 4.480 44.800 4.760 ;
      LAYER met1 ;
        RECT 44.800 4.480 46.480 4.760 ;
      LAYER met1 ;
        RECT 0.000 4.200 42.840 4.480 ;
      LAYER met1 ;
        RECT 42.840 4.200 46.480 4.480 ;
      LAYER met1 ;
        RECT 46.480 4.200 52.360 5.040 ;
      LAYER met1 ;
        RECT 52.360 4.760 53.200 5.600 ;
      LAYER met1 ;
        RECT 53.200 4.760 92.400 5.600 ;
      LAYER met1 ;
        RECT 52.360 4.480 54.600 4.760 ;
      LAYER met1 ;
        RECT 54.600 4.480 92.400 4.760 ;
      LAYER met1 ;
        RECT 52.360 4.200 56.560 4.480 ;
      LAYER met1 ;
        RECT 56.560 4.200 92.400 4.480 ;
        RECT 0.000 3.920 42.560 4.200 ;
      LAYER met1 ;
        RECT 42.560 3.920 44.800 4.200 ;
      LAYER met1 ;
        RECT 44.800 3.920 45.640 4.200 ;
      LAYER met1 ;
        RECT 45.640 3.920 46.480 4.200 ;
      LAYER met1 ;
        RECT 46.480 3.920 47.880 4.200 ;
      LAYER met1 ;
        RECT 47.880 3.920 48.160 4.200 ;
      LAYER met1 ;
        RECT 0.000 3.640 42.280 3.920 ;
      LAYER met1 ;
        RECT 42.280 3.640 42.840 3.920 ;
      LAYER met1 ;
        RECT 42.840 3.640 45.640 3.920 ;
      LAYER met1 ;
        RECT 45.640 3.640 46.760 3.920 ;
      LAYER met1 ;
        RECT 46.760 3.640 47.600 3.920 ;
      LAYER met1 ;
        RECT 47.600 3.640 48.160 3.920 ;
      LAYER met1 ;
        RECT 48.160 3.640 49.280 4.200 ;
      LAYER met1 ;
        RECT 49.280 3.920 49.560 4.200 ;
      LAYER met1 ;
        RECT 49.560 3.920 50.960 4.200 ;
      LAYER met1 ;
        RECT 50.960 3.920 51.240 4.200 ;
      LAYER met1 ;
        RECT 51.240 3.920 52.360 4.200 ;
      LAYER met1 ;
        RECT 52.360 3.920 53.200 4.200 ;
      LAYER met1 ;
        RECT 53.200 3.920 54.600 4.200 ;
      LAYER met1 ;
        RECT 54.600 3.920 56.840 4.200 ;
      LAYER met1 ;
        RECT 56.840 3.920 92.400 4.200 ;
      LAYER met1 ;
        RECT 49.280 3.640 49.840 3.920 ;
      LAYER met1 ;
        RECT 0.000 3.360 42.000 3.640 ;
      LAYER met1 ;
        RECT 42.000 3.360 42.560 3.640 ;
      LAYER met1 ;
        RECT 0.000 3.080 41.720 3.360 ;
      LAYER met1 ;
        RECT 41.720 3.080 42.560 3.360 ;
      LAYER met1 ;
        RECT 42.560 3.080 45.360 3.640 ;
        RECT 0.000 2.520 41.440 3.080 ;
      LAYER met1 ;
        RECT 41.440 2.800 42.280 3.080 ;
      LAYER met1 ;
        RECT 42.280 2.800 45.360 3.080 ;
      LAYER met1 ;
        RECT 45.360 2.800 45.920 3.640 ;
      LAYER met1 ;
        RECT 45.920 3.360 46.200 3.640 ;
      LAYER met1 ;
        RECT 46.200 3.360 46.760 3.640 ;
      LAYER met1 ;
        RECT 46.760 3.360 47.320 3.640 ;
      LAYER met1 ;
        RECT 47.320 3.360 48.160 3.640 ;
      LAYER met1 ;
        RECT 48.160 3.360 49.000 3.640 ;
      LAYER met1 ;
        RECT 49.000 3.360 49.840 3.640 ;
      LAYER met1 ;
        RECT 49.840 3.360 50.960 3.920 ;
      LAYER met1 ;
        RECT 50.960 3.640 51.520 3.920 ;
      LAYER met1 ;
        RECT 51.520 3.640 52.640 3.920 ;
      LAYER met1 ;
        RECT 52.640 3.640 53.200 3.920 ;
      LAYER met1 ;
        RECT 53.200 3.640 56.280 3.920 ;
      LAYER met1 ;
        RECT 56.280 3.640 57.120 3.920 ;
      LAYER met1 ;
        RECT 57.120 3.640 92.400 3.920 ;
      LAYER met1 ;
        RECT 50.960 3.360 51.800 3.640 ;
      LAYER met1 ;
        RECT 51.800 3.360 52.640 3.640 ;
      LAYER met1 ;
        RECT 52.640 3.360 53.480 3.640 ;
      LAYER met1 ;
        RECT 53.480 3.360 56.560 3.640 ;
      LAYER met1 ;
        RECT 56.560 3.360 57.400 3.640 ;
      LAYER met1 ;
        RECT 57.400 3.360 92.400 3.640 ;
        RECT 45.920 2.800 46.480 3.360 ;
      LAYER met1 ;
        RECT 46.480 2.800 47.600 3.360 ;
      LAYER met1 ;
        RECT 47.600 3.080 47.880 3.360 ;
      LAYER met1 ;
        RECT 47.880 3.080 48.440 3.360 ;
      LAYER met1 ;
        RECT 48.440 3.080 49.000 3.360 ;
      LAYER met1 ;
        RECT 49.000 3.080 49.280 3.360 ;
      LAYER met1 ;
        RECT 49.280 3.080 49.560 3.360 ;
      LAYER met1 ;
        RECT 49.560 3.080 50.120 3.360 ;
      LAYER met1 ;
        RECT 47.600 2.800 48.160 3.080 ;
      LAYER met1 ;
        RECT 48.160 2.800 48.440 3.080 ;
      LAYER met1 ;
        RECT 48.440 2.800 48.720 3.080 ;
      LAYER met1 ;
        RECT 48.720 2.800 49.280 3.080 ;
      LAYER met1 ;
        RECT 49.280 2.800 49.840 3.080 ;
      LAYER met1 ;
        RECT 49.840 2.800 50.120 3.080 ;
      LAYER met1 ;
        RECT 50.120 2.800 50.680 3.360 ;
      LAYER met1 ;
        RECT 50.680 3.080 51.240 3.360 ;
      LAYER met1 ;
        RECT 51.240 3.080 51.520 3.360 ;
      LAYER met1 ;
        RECT 51.520 3.080 51.800 3.360 ;
      LAYER met1 ;
        RECT 51.800 3.080 52.360 3.360 ;
      LAYER met1 ;
        RECT 52.360 3.080 53.480 3.360 ;
      LAYER met1 ;
        RECT 53.480 3.080 56.840 3.360 ;
      LAYER met1 ;
        RECT 56.840 3.080 57.680 3.360 ;
        RECT 50.680 2.800 50.960 3.080 ;
      LAYER met1 ;
        RECT 50.960 2.800 51.520 3.080 ;
      LAYER met1 ;
        RECT 51.520 2.800 52.080 3.080 ;
      LAYER met1 ;
        RECT 52.080 2.800 52.360 3.080 ;
      LAYER met1 ;
        RECT 52.360 2.800 53.760 3.080 ;
      LAYER met1 ;
        RECT 53.760 2.800 57.120 3.080 ;
      LAYER met1 ;
        RECT 57.120 2.800 57.680 3.080 ;
      LAYER met1 ;
        RECT 57.680 2.800 92.400 3.360 ;
      LAYER met1 ;
        RECT 41.440 2.520 42.000 2.800 ;
      LAYER met1 ;
        RECT 42.000 2.520 45.360 2.800 ;
      LAYER met1 ;
        RECT 45.360 2.520 46.200 2.800 ;
      LAYER met1 ;
        RECT 46.200 2.520 46.760 2.800 ;
      LAYER met1 ;
        RECT 46.760 2.520 47.320 2.800 ;
      LAYER met1 ;
        RECT 0.000 2.240 41.160 2.520 ;
      LAYER met1 ;
        RECT 41.160 2.240 41.720 2.520 ;
      LAYER met1 ;
        RECT 41.720 2.240 45.080 2.520 ;
      LAYER met1 ;
        RECT 45.080 2.240 47.320 2.520 ;
      LAYER met1 ;
        RECT 47.320 2.240 48.160 2.800 ;
      LAYER met1 ;
        RECT 48.160 2.240 49.000 2.800 ;
      LAYER met1 ;
        RECT 49.000 2.520 49.840 2.800 ;
      LAYER met1 ;
        RECT 49.840 2.520 50.960 2.800 ;
      LAYER met1 ;
        RECT 50.960 2.520 51.800 2.800 ;
      LAYER met1 ;
        RECT 51.800 2.520 54.040 2.800 ;
      LAYER met1 ;
        RECT 54.040 2.520 57.400 2.800 ;
      LAYER met1 ;
        RECT 57.400 2.520 57.960 2.800 ;
      LAYER met1 ;
        RECT 57.960 2.520 92.400 2.800 ;
        RECT 49.000 2.240 50.120 2.520 ;
      LAYER met1 ;
        RECT 50.120 2.240 50.680 2.520 ;
      LAYER met1 ;
        RECT 50.680 2.240 51.800 2.520 ;
      LAYER met1 ;
        RECT 51.800 2.240 53.480 2.520 ;
      LAYER met1 ;
        RECT 53.480 2.240 53.760 2.520 ;
      LAYER met1 ;
        RECT 53.760 2.240 54.320 2.520 ;
      LAYER met1 ;
        RECT 54.320 2.240 57.680 2.520 ;
      LAYER met1 ;
        RECT 57.680 2.240 58.240 2.520 ;
      LAYER met1 ;
        RECT 58.240 2.240 92.400 2.520 ;
        RECT 0.000 1.960 40.880 2.240 ;
      LAYER met1 ;
        RECT 40.880 1.960 41.440 2.240 ;
      LAYER met1 ;
        RECT 41.440 1.960 44.800 2.240 ;
      LAYER met1 ;
        RECT 44.800 1.960 45.360 2.240 ;
      LAYER met1 ;
        RECT 45.360 1.960 45.920 2.240 ;
      LAYER met1 ;
        RECT 45.920 1.960 53.480 2.240 ;
      LAYER met1 ;
        RECT 53.480 1.960 54.040 2.240 ;
      LAYER met1 ;
        RECT 54.040 1.960 54.600 2.240 ;
      LAYER met1 ;
        RECT 54.600 1.960 57.960 2.240 ;
      LAYER met1 ;
        RECT 57.960 1.960 58.520 2.240 ;
      LAYER met1 ;
        RECT 58.520 1.960 92.400 2.240 ;
        RECT 0.000 1.680 40.600 1.960 ;
      LAYER met1 ;
        RECT 40.600 1.680 41.160 1.960 ;
      LAYER met1 ;
        RECT 41.160 1.680 44.520 1.960 ;
      LAYER met1 ;
        RECT 44.520 1.680 45.080 1.960 ;
      LAYER met1 ;
        RECT 45.080 1.680 45.920 1.960 ;
      LAYER met1 ;
        RECT 45.920 1.680 53.200 1.960 ;
      LAYER met1 ;
        RECT 53.200 1.680 54.320 1.960 ;
      LAYER met1 ;
        RECT 54.320 1.680 54.880 1.960 ;
      LAYER met1 ;
        RECT 54.880 1.680 58.240 1.960 ;
      LAYER met1 ;
        RECT 58.240 1.680 58.800 1.960 ;
      LAYER met1 ;
        RECT 58.800 1.680 92.400 1.960 ;
        RECT 0.000 1.400 40.320 1.680 ;
      LAYER met1 ;
        RECT 40.320 1.400 40.880 1.680 ;
      LAYER met1 ;
        RECT 40.880 1.400 43.400 1.680 ;
      LAYER met1 ;
        RECT 43.400 1.400 44.800 1.680 ;
      LAYER met1 ;
        RECT 44.800 1.400 45.920 1.680 ;
      LAYER met1 ;
        RECT 45.920 1.400 46.760 1.680 ;
      LAYER met1 ;
        RECT 46.760 1.400 47.320 1.680 ;
      LAYER met1 ;
        RECT 47.320 1.400 47.880 1.680 ;
      LAYER met1 ;
        RECT 0.000 1.120 40.040 1.400 ;
      LAYER met1 ;
        RECT 40.040 1.120 40.600 1.400 ;
      LAYER met1 ;
        RECT 40.600 1.120 41.160 1.400 ;
      LAYER met1 ;
        RECT 41.160 1.120 44.520 1.400 ;
      LAYER met1 ;
        RECT 44.520 1.120 45.920 1.400 ;
      LAYER met1 ;
        RECT 45.920 1.120 47.880 1.400 ;
      LAYER met1 ;
        RECT 47.880 1.120 50.680 1.680 ;
      LAYER met1 ;
        RECT 50.680 1.400 51.520 1.680 ;
      LAYER met1 ;
        RECT 51.520 1.400 52.080 1.680 ;
      LAYER met1 ;
        RECT 52.080 1.400 52.920 1.680 ;
      LAYER met1 ;
        RECT 52.920 1.400 54.600 1.680 ;
      LAYER met1 ;
        RECT 54.600 1.400 56.000 1.680 ;
      LAYER met1 ;
        RECT 56.000 1.400 58.520 1.680 ;
      LAYER met1 ;
        RECT 58.520 1.400 59.080 1.680 ;
      LAYER met1 ;
        RECT 59.080 1.400 92.400 1.680 ;
      LAYER met1 ;
        RECT 50.680 1.120 52.640 1.400 ;
      LAYER met1 ;
        RECT 52.640 1.120 54.880 1.400 ;
      LAYER met1 ;
        RECT 54.880 1.120 57.960 1.400 ;
      LAYER met1 ;
        RECT 57.960 1.120 58.800 1.400 ;
      LAYER met1 ;
        RECT 58.800 1.120 59.360 1.400 ;
      LAYER met1 ;
        RECT 59.360 1.120 92.400 1.400 ;
        RECT 0.000 0.560 39.760 1.120 ;
      LAYER met1 ;
        RECT 39.760 0.840 43.400 1.120 ;
      LAYER met1 ;
        RECT 43.400 0.840 46.200 1.120 ;
      LAYER met1 ;
        RECT 46.200 0.840 47.600 1.120 ;
      LAYER met1 ;
        RECT 47.600 0.840 50.960 1.120 ;
      LAYER met1 ;
        RECT 50.960 0.840 52.640 1.120 ;
      LAYER met1 ;
        RECT 52.640 0.840 56.000 1.120 ;
      LAYER met1 ;
        RECT 56.000 0.840 59.640 1.120 ;
        RECT 39.760 0.560 41.160 0.840 ;
      LAYER met1 ;
        RECT 41.160 0.560 51.240 0.840 ;
      LAYER met1 ;
        RECT 51.240 0.560 52.080 0.840 ;
      LAYER met1 ;
        RECT 52.080 0.560 57.960 0.840 ;
      LAYER met1 ;
        RECT 57.960 0.560 59.640 0.840 ;
      LAYER met1 ;
        RECT 59.640 0.560 92.400 1.120 ;
        RECT 0.000 0.000 92.400 0.560 ;
      LAYER met2 ;
        RECT 0.000 28.840 92.400 29.400 ;
        RECT 0.000 28.560 44.240 28.840 ;
      LAYER met2 ;
        RECT 44.240 28.560 45.080 28.840 ;
      LAYER met2 ;
        RECT 45.080 28.560 92.400 28.840 ;
        RECT 0.000 26.040 43.960 28.560 ;
      LAYER met2 ;
        RECT 43.960 28.280 45.920 28.560 ;
      LAYER met2 ;
        RECT 45.920 28.280 92.400 28.560 ;
      LAYER met2 ;
        RECT 43.960 26.040 44.520 28.280 ;
      LAYER met2 ;
        RECT 44.520 28.000 45.080 28.280 ;
      LAYER met2 ;
        RECT 45.080 28.000 46.480 28.280 ;
      LAYER met2 ;
        RECT 46.480 28.000 92.400 28.280 ;
        RECT 44.520 27.720 45.920 28.000 ;
      LAYER met2 ;
        RECT 45.920 27.720 47.320 28.000 ;
      LAYER met2 ;
        RECT 47.320 27.720 92.400 28.000 ;
        RECT 44.520 27.440 46.480 27.720 ;
      LAYER met2 ;
        RECT 46.480 27.440 47.880 27.720 ;
      LAYER met2 ;
        RECT 47.880 27.440 53.760 27.720 ;
      LAYER met2 ;
        RECT 53.760 27.440 56.280 27.720 ;
      LAYER met2 ;
        RECT 56.280 27.440 92.400 27.720 ;
        RECT 44.520 27.160 47.320 27.440 ;
      LAYER met2 ;
        RECT 47.320 27.160 48.440 27.440 ;
      LAYER met2 ;
        RECT 48.440 27.160 52.360 27.440 ;
      LAYER met2 ;
        RECT 52.360 27.160 56.560 27.440 ;
      LAYER met2 ;
        RECT 44.520 26.880 47.880 27.160 ;
      LAYER met2 ;
        RECT 47.880 26.880 49.000 27.160 ;
      LAYER met2 ;
        RECT 49.000 26.880 49.280 27.160 ;
      LAYER met2 ;
        RECT 49.280 26.880 50.400 27.160 ;
      LAYER met2 ;
        RECT 50.400 26.880 51.240 27.160 ;
      LAYER met2 ;
        RECT 51.240 26.880 53.760 27.160 ;
      LAYER met2 ;
        RECT 53.760 26.880 56.000 27.160 ;
        RECT 44.520 26.600 48.440 26.880 ;
      LAYER met2 ;
        RECT 48.440 26.600 52.360 26.880 ;
      LAYER met2 ;
        RECT 52.360 26.600 56.000 26.880 ;
        RECT 44.520 26.320 48.720 26.600 ;
      LAYER met2 ;
        RECT 48.720 26.320 49.560 26.600 ;
      LAYER met2 ;
        RECT 49.560 26.320 50.120 26.600 ;
      LAYER met2 ;
        RECT 50.120 26.320 51.240 26.600 ;
      LAYER met2 ;
        RECT 51.240 26.320 56.000 26.600 ;
        RECT 44.520 26.040 48.440 26.320 ;
      LAYER met2 ;
        RECT 48.440 26.040 50.960 26.320 ;
      LAYER met2 ;
        RECT 50.960 26.040 56.000 26.320 ;
        RECT 0.000 25.760 43.400 26.040 ;
      LAYER met2 ;
        RECT 43.400 25.760 44.520 26.040 ;
      LAYER met2 ;
        RECT 44.520 25.760 47.040 26.040 ;
      LAYER met2 ;
        RECT 47.040 25.760 52.080 26.040 ;
      LAYER met2 ;
        RECT 52.080 25.760 56.000 26.040 ;
        RECT 0.000 25.480 42.840 25.760 ;
      LAYER met2 ;
        RECT 42.840 25.480 43.960 25.760 ;
      LAYER met2 ;
        RECT 43.960 25.480 44.240 25.760 ;
        RECT 0.000 25.200 5.880 25.480 ;
      LAYER met2 ;
        RECT 5.880 25.200 9.800 25.480 ;
      LAYER met2 ;
        RECT 9.800 25.200 23.240 25.480 ;
      LAYER met2 ;
        RECT 23.240 25.200 27.160 25.480 ;
      LAYER met2 ;
        RECT 27.160 25.200 42.280 25.480 ;
      LAYER met2 ;
        RECT 42.280 25.200 43.400 25.480 ;
      LAYER met2 ;
        RECT 43.400 25.200 44.240 25.480 ;
      LAYER met2 ;
        RECT 44.240 25.200 44.800 25.760 ;
      LAYER met2 ;
        RECT 44.800 25.480 45.920 25.760 ;
      LAYER met2 ;
        RECT 45.920 25.480 48.440 25.760 ;
      LAYER met2 ;
        RECT 48.440 25.480 50.960 25.760 ;
      LAYER met2 ;
        RECT 50.960 25.480 52.640 25.760 ;
      LAYER met2 ;
        RECT 52.640 25.480 56.000 25.760 ;
        RECT 44.800 25.200 45.080 25.480 ;
      LAYER met2 ;
        RECT 45.080 25.200 47.040 25.480 ;
      LAYER met2 ;
        RECT 47.040 25.200 52.080 25.480 ;
      LAYER met2 ;
        RECT 52.080 25.200 53.200 25.480 ;
      LAYER met2 ;
        RECT 53.200 25.200 56.000 25.480 ;
      LAYER met2 ;
        RECT 56.000 25.200 56.560 27.160 ;
      LAYER met2 ;
        RECT 56.560 25.200 92.400 27.440 ;
        RECT 0.000 24.920 5.040 25.200 ;
      LAYER met2 ;
        RECT 5.040 24.920 10.360 25.200 ;
      LAYER met2 ;
        RECT 10.360 24.920 22.400 25.200 ;
      LAYER met2 ;
        RECT 22.400 24.920 28.000 25.200 ;
      LAYER met2 ;
        RECT 28.000 24.920 42.000 25.200 ;
      LAYER met2 ;
        RECT 42.000 24.920 42.840 25.200 ;
      LAYER met2 ;
        RECT 42.840 24.920 44.240 25.200 ;
      LAYER met2 ;
        RECT 44.240 24.920 45.920 25.200 ;
      LAYER met2 ;
        RECT 45.920 24.920 52.640 25.200 ;
      LAYER met2 ;
        RECT 52.640 24.920 53.760 25.200 ;
      LAYER met2 ;
        RECT 53.760 24.920 55.720 25.200 ;
        RECT 0.000 24.640 4.480 24.920 ;
      LAYER met2 ;
        RECT 4.480 24.640 10.920 24.920 ;
      LAYER met2 ;
        RECT 10.920 24.640 21.840 24.920 ;
      LAYER met2 ;
        RECT 21.840 24.640 28.560 24.920 ;
      LAYER met2 ;
        RECT 28.560 24.640 41.720 24.920 ;
      LAYER met2 ;
        RECT 41.720 24.640 42.560 24.920 ;
      LAYER met2 ;
        RECT 42.560 24.640 43.960 24.920 ;
      LAYER met2 ;
        RECT 43.960 24.640 45.080 24.920 ;
      LAYER met2 ;
        RECT 45.080 24.640 53.200 24.920 ;
      LAYER met2 ;
        RECT 53.200 24.640 54.040 24.920 ;
      LAYER met2 ;
        RECT 54.040 24.640 55.720 24.920 ;
      LAYER met2 ;
        RECT 55.720 24.640 56.280 25.200 ;
      LAYER met2 ;
        RECT 56.280 24.640 92.400 25.200 ;
        RECT 0.000 24.360 3.920 24.640 ;
      LAYER met2 ;
        RECT 3.920 24.360 11.480 24.640 ;
      LAYER met2 ;
        RECT 11.480 24.360 21.280 24.640 ;
      LAYER met2 ;
        RECT 21.280 24.360 29.120 24.640 ;
      LAYER met2 ;
        RECT 29.120 24.360 41.720 24.640 ;
      LAYER met2 ;
        RECT 41.720 24.360 43.120 24.640 ;
      LAYER met2 ;
        RECT 43.120 24.360 43.680 24.640 ;
      LAYER met2 ;
        RECT 43.680 24.360 44.520 24.640 ;
      LAYER met2 ;
        RECT 44.520 24.360 53.480 24.640 ;
      LAYER met2 ;
        RECT 53.480 24.360 54.320 24.640 ;
      LAYER met2 ;
        RECT 54.320 24.360 55.440 24.640 ;
      LAYER met2 ;
        RECT 55.440 24.360 56.560 24.640 ;
      LAYER met2 ;
        RECT 56.560 24.360 92.400 24.640 ;
        RECT 0.000 24.080 3.360 24.360 ;
      LAYER met2 ;
        RECT 3.360 24.080 6.160 24.360 ;
      LAYER met2 ;
        RECT 6.160 24.080 9.240 24.360 ;
      LAYER met2 ;
        RECT 9.240 24.080 12.040 24.360 ;
      LAYER met2 ;
        RECT 12.040 24.080 21.000 24.360 ;
      LAYER met2 ;
        RECT 21.000 24.080 23.800 24.360 ;
      LAYER met2 ;
        RECT 23.800 24.080 26.600 24.360 ;
      LAYER met2 ;
        RECT 26.600 24.080 29.400 24.360 ;
      LAYER met2 ;
        RECT 29.400 24.080 42.560 24.360 ;
      LAYER met2 ;
        RECT 42.560 24.080 44.240 24.360 ;
      LAYER met2 ;
        RECT 44.240 24.080 54.040 24.360 ;
      LAYER met2 ;
        RECT 54.040 24.080 54.600 24.360 ;
      LAYER met2 ;
        RECT 54.600 24.080 55.440 24.360 ;
      LAYER met2 ;
        RECT 55.440 24.080 56.840 24.360 ;
      LAYER met2 ;
        RECT 56.840 24.080 92.400 24.360 ;
        RECT 0.000 23.800 3.080 24.080 ;
      LAYER met2 ;
        RECT 3.080 23.800 5.320 24.080 ;
      LAYER met2 ;
        RECT 5.320 23.800 10.080 24.080 ;
      LAYER met2 ;
        RECT 10.080 23.800 12.320 24.080 ;
      LAYER met2 ;
        RECT 12.320 23.800 20.720 24.080 ;
      LAYER met2 ;
        RECT 20.720 23.800 22.960 24.080 ;
      LAYER met2 ;
        RECT 22.960 23.800 27.440 24.080 ;
      LAYER met2 ;
        RECT 27.440 23.800 29.680 24.080 ;
      LAYER met2 ;
        RECT 29.680 23.800 42.840 24.080 ;
      LAYER met2 ;
        RECT 42.840 23.800 43.680 24.080 ;
      LAYER met2 ;
        RECT 43.680 23.800 54.320 24.080 ;
      LAYER met2 ;
        RECT 54.320 23.800 54.880 24.080 ;
      LAYER met2 ;
        RECT 54.880 23.800 55.160 24.080 ;
      LAYER met2 ;
        RECT 55.160 23.800 56.000 24.080 ;
      LAYER met2 ;
        RECT 56.000 23.800 56.280 24.080 ;
      LAYER met2 ;
        RECT 56.280 23.800 57.120 24.080 ;
      LAYER met2 ;
        RECT 57.120 23.800 92.400 24.080 ;
        RECT 0.000 23.520 2.800 23.800 ;
      LAYER met2 ;
        RECT 2.800 23.520 4.760 23.800 ;
      LAYER met2 ;
        RECT 4.760 23.520 10.640 23.800 ;
      LAYER met2 ;
        RECT 10.640 23.520 12.600 23.800 ;
      LAYER met2 ;
        RECT 12.600 23.520 20.440 23.800 ;
      LAYER met2 ;
        RECT 20.440 23.520 22.400 23.800 ;
      LAYER met2 ;
        RECT 22.400 23.520 28.000 23.800 ;
      LAYER met2 ;
        RECT 28.000 23.520 29.960 23.800 ;
      LAYER met2 ;
        RECT 29.960 23.520 42.560 23.800 ;
      LAYER met2 ;
        RECT 42.560 23.520 43.400 23.800 ;
      LAYER met2 ;
        RECT 43.400 23.520 54.600 23.800 ;
      LAYER met2 ;
        RECT 54.600 23.520 55.720 23.800 ;
      LAYER met2 ;
        RECT 55.720 23.520 56.560 23.800 ;
      LAYER met2 ;
        RECT 56.560 23.520 57.400 23.800 ;
      LAYER met2 ;
        RECT 57.400 23.520 92.400 23.800 ;
        RECT 0.000 23.240 2.520 23.520 ;
      LAYER met2 ;
        RECT 2.520 23.240 4.480 23.520 ;
      LAYER met2 ;
        RECT 4.480 23.240 10.920 23.520 ;
      LAYER met2 ;
        RECT 10.920 23.240 12.880 23.520 ;
      LAYER met2 ;
        RECT 12.880 23.240 20.160 23.520 ;
      LAYER met2 ;
        RECT 20.160 23.240 21.840 23.520 ;
      LAYER met2 ;
        RECT 21.840 23.240 28.560 23.520 ;
      LAYER met2 ;
        RECT 28.560 23.240 30.240 23.520 ;
      LAYER met2 ;
        RECT 30.240 23.240 42.560 23.520 ;
        RECT 0.000 22.960 2.240 23.240 ;
      LAYER met2 ;
        RECT 2.240 22.960 3.920 23.240 ;
      LAYER met2 ;
        RECT 3.920 22.960 11.480 23.240 ;
      LAYER met2 ;
        RECT 11.480 22.960 13.160 23.240 ;
      LAYER met2 ;
        RECT 13.160 22.960 19.880 23.240 ;
      LAYER met2 ;
        RECT 19.880 22.960 21.560 23.240 ;
      LAYER met2 ;
        RECT 21.560 22.960 28.840 23.240 ;
      LAYER met2 ;
        RECT 28.840 22.960 30.520 23.240 ;
      LAYER met2 ;
        RECT 30.520 22.960 42.560 23.240 ;
      LAYER met2 ;
        RECT 42.560 22.960 43.120 23.520 ;
      LAYER met2 ;
        RECT 43.120 22.960 54.880 23.520 ;
      LAYER met2 ;
        RECT 54.880 22.960 55.440 23.520 ;
      LAYER met2 ;
        RECT 55.440 23.240 56.840 23.520 ;
      LAYER met2 ;
        RECT 56.840 23.240 57.680 23.520 ;
      LAYER met2 ;
        RECT 57.680 23.240 92.400 23.520 ;
        RECT 55.440 22.960 57.120 23.240 ;
      LAYER met2 ;
        RECT 57.120 22.960 57.960 23.240 ;
      LAYER met2 ;
        RECT 57.960 22.960 92.400 23.240 ;
        RECT 0.000 22.680 1.960 22.960 ;
      LAYER met2 ;
        RECT 1.960 22.680 3.640 22.960 ;
      LAYER met2 ;
        RECT 3.640 22.680 11.760 22.960 ;
      LAYER met2 ;
        RECT 11.760 22.680 13.440 22.960 ;
      LAYER met2 ;
        RECT 13.440 22.680 19.600 22.960 ;
      LAYER met2 ;
        RECT 19.600 22.680 21.280 22.960 ;
      LAYER met2 ;
        RECT 21.280 22.680 29.120 22.960 ;
      LAYER met2 ;
        RECT 29.120 22.680 30.800 22.960 ;
      LAYER met2 ;
        RECT 30.800 22.680 42.280 22.960 ;
        RECT 0.000 22.120 1.680 22.680 ;
      LAYER met2 ;
        RECT 1.680 22.120 8.960 22.680 ;
      LAYER met2 ;
        RECT 8.960 22.400 12.040 22.680 ;
      LAYER met2 ;
        RECT 12.040 22.400 13.440 22.680 ;
      LAYER met2 ;
        RECT 13.440 22.400 19.320 22.680 ;
      LAYER met2 ;
        RECT 19.320 22.400 21.000 22.680 ;
      LAYER met2 ;
        RECT 21.000 22.400 24.920 22.680 ;
      LAYER met2 ;
        RECT 24.920 22.400 26.040 22.680 ;
      LAYER met2 ;
        RECT 26.040 22.400 29.400 22.680 ;
      LAYER met2 ;
        RECT 29.400 22.400 31.080 22.680 ;
      LAYER met2 ;
        RECT 31.080 22.400 42.280 22.680 ;
        RECT 0.000 21.560 1.400 22.120 ;
      LAYER met2 ;
        RECT 1.400 21.560 8.960 22.120 ;
      LAYER met2 ;
        RECT 8.960 21.840 12.320 22.400 ;
      LAYER met2 ;
        RECT 12.320 22.120 13.720 22.400 ;
      LAYER met2 ;
        RECT 13.720 22.120 19.320 22.400 ;
      LAYER met2 ;
        RECT 19.320 22.120 20.720 22.400 ;
      LAYER met2 ;
        RECT 20.720 22.120 24.080 22.400 ;
      LAYER met2 ;
        RECT 24.080 22.120 26.880 22.400 ;
      LAYER met2 ;
        RECT 26.880 22.120 29.680 22.400 ;
      LAYER met2 ;
        RECT 29.680 22.120 31.360 22.400 ;
      LAYER met2 ;
        RECT 31.360 22.120 42.280 22.400 ;
      LAYER met2 ;
        RECT 42.280 22.120 42.840 22.960 ;
      LAYER met2 ;
        RECT 42.840 22.680 55.160 22.960 ;
      LAYER met2 ;
        RECT 55.160 22.680 55.720 22.960 ;
      LAYER met2 ;
        RECT 55.720 22.680 57.120 22.960 ;
      LAYER met2 ;
        RECT 57.120 22.680 58.240 22.960 ;
      LAYER met2 ;
        RECT 42.840 22.400 55.440 22.680 ;
        RECT 42.840 22.120 47.040 22.400 ;
      LAYER met2 ;
        RECT 47.040 22.120 47.320 22.400 ;
      LAYER met2 ;
        RECT 47.320 22.120 55.440 22.400 ;
      LAYER met2 ;
        RECT 55.440 22.120 56.000 22.680 ;
      LAYER met2 ;
        RECT 56.000 22.400 56.560 22.680 ;
      LAYER met2 ;
        RECT 56.560 22.400 58.240 22.680 ;
      LAYER met2 ;
        RECT 58.240 22.400 92.400 22.960 ;
        RECT 56.000 22.120 56.280 22.400 ;
      LAYER met2 ;
        RECT 56.280 22.120 57.400 22.400 ;
      LAYER met2 ;
        RECT 57.400 22.120 71.960 22.400 ;
      LAYER met2 ;
        RECT 71.960 22.120 72.800 22.400 ;
      LAYER met2 ;
        RECT 72.800 22.120 92.400 22.400 ;
      LAYER met2 ;
        RECT 12.320 21.840 14.000 22.120 ;
      LAYER met2 ;
        RECT 14.000 21.840 19.040 22.120 ;
      LAYER met2 ;
        RECT 19.040 21.840 20.440 22.120 ;
      LAYER met2 ;
        RECT 20.440 21.840 23.520 22.120 ;
      LAYER met2 ;
        RECT 23.520 21.840 27.160 22.120 ;
      LAYER met2 ;
        RECT 27.160 21.840 29.960 22.120 ;
      LAYER met2 ;
        RECT 29.960 21.840 31.360 22.120 ;
      LAYER met2 ;
        RECT 31.360 21.840 42.000 22.120 ;
      LAYER met2 ;
        RECT 42.000 21.840 42.840 22.120 ;
      LAYER met2 ;
        RECT 42.840 21.840 44.520 22.120 ;
      LAYER met2 ;
        RECT 44.520 21.840 44.800 22.120 ;
      LAYER met2 ;
        RECT 44.800 21.840 45.920 22.120 ;
      LAYER met2 ;
        RECT 45.920 21.840 46.200 22.120 ;
      LAYER met2 ;
        RECT 8.960 21.560 12.600 21.840 ;
      LAYER met2 ;
        RECT 12.600 21.560 14.000 21.840 ;
      LAYER met2 ;
        RECT 14.000 21.560 18.760 21.840 ;
        RECT 0.000 20.720 1.120 21.560 ;
      LAYER met2 ;
        RECT 1.120 20.720 8.960 21.560 ;
      LAYER met2 ;
        RECT 8.960 21.000 12.880 21.560 ;
      LAYER met2 ;
        RECT 12.880 21.000 14.280 21.560 ;
      LAYER met2 ;
        RECT 14.280 21.000 18.760 21.560 ;
      LAYER met2 ;
        RECT 18.760 21.280 20.160 21.840 ;
      LAYER met2 ;
        RECT 20.160 21.560 23.240 21.840 ;
      LAYER met2 ;
        RECT 23.240 21.560 27.440 21.840 ;
      LAYER met2 ;
        RECT 27.440 21.560 30.240 21.840 ;
        RECT 20.160 21.280 22.960 21.560 ;
      LAYER met2 ;
        RECT 22.960 21.280 27.720 21.560 ;
      LAYER met2 ;
        RECT 27.720 21.280 30.240 21.560 ;
      LAYER met2 ;
        RECT 30.240 21.280 31.640 21.840 ;
      LAYER met2 ;
        RECT 31.640 21.560 42.000 21.840 ;
      LAYER met2 ;
        RECT 42.000 21.560 42.560 21.840 ;
      LAYER met2 ;
        RECT 31.640 21.280 41.720 21.560 ;
      LAYER met2 ;
        RECT 41.720 21.280 42.560 21.560 ;
      LAYER met2 ;
        RECT 42.560 21.280 44.240 21.840 ;
      LAYER met2 ;
        RECT 44.240 21.280 44.800 21.840 ;
      LAYER met2 ;
        RECT 44.800 21.560 45.640 21.840 ;
      LAYER met2 ;
        RECT 45.640 21.560 46.200 21.840 ;
      LAYER met2 ;
        RECT 46.200 21.560 46.760 22.120 ;
      LAYER met2 ;
        RECT 46.760 21.560 47.320 22.120 ;
      LAYER met2 ;
        RECT 47.320 21.840 49.280 22.120 ;
      LAYER met2 ;
        RECT 49.280 21.840 49.840 22.120 ;
      LAYER met2 ;
        RECT 49.840 21.840 55.720 22.120 ;
      LAYER met2 ;
        RECT 55.720 21.840 56.840 22.120 ;
      LAYER met2 ;
        RECT 56.840 21.840 71.680 22.120 ;
      LAYER met2 ;
        RECT 71.680 21.840 72.800 22.120 ;
      LAYER met2 ;
        RECT 72.800 21.840 79.520 22.120 ;
      LAYER met2 ;
        RECT 79.520 21.840 80.080 22.120 ;
      LAYER met2 ;
        RECT 80.080 21.840 91.000 22.120 ;
      LAYER met2 ;
        RECT 91.000 21.840 91.560 22.120 ;
      LAYER met2 ;
        RECT 91.560 21.840 92.400 22.120 ;
        RECT 47.320 21.560 49.000 21.840 ;
      LAYER met2 ;
        RECT 49.000 21.560 49.840 21.840 ;
      LAYER met2 ;
        RECT 49.840 21.560 50.680 21.840 ;
      LAYER met2 ;
        RECT 50.680 21.560 50.960 21.840 ;
      LAYER met2 ;
        RECT 50.960 21.560 52.080 21.840 ;
      LAYER met2 ;
        RECT 52.080 21.560 52.360 21.840 ;
      LAYER met2 ;
        RECT 52.360 21.560 55.720 21.840 ;
      LAYER met2 ;
        RECT 18.760 21.000 19.880 21.280 ;
      LAYER met2 ;
        RECT 19.880 21.000 22.960 21.280 ;
      LAYER met2 ;
        RECT 22.960 21.000 28.000 21.280 ;
      LAYER met2 ;
        RECT 8.960 20.720 13.160 21.000 ;
      LAYER met2 ;
        RECT 13.160 20.720 14.280 21.000 ;
      LAYER met2 ;
        RECT 14.280 20.720 18.480 21.000 ;
      LAYER met2 ;
        RECT 18.480 20.720 19.880 21.000 ;
      LAYER met2 ;
        RECT 19.880 20.720 22.680 21.000 ;
      LAYER met2 ;
        RECT 22.680 20.720 24.920 21.000 ;
      LAYER met2 ;
        RECT 24.920 20.720 26.040 21.000 ;
      LAYER met2 ;
        RECT 26.040 20.720 28.000 21.000 ;
      LAYER met2 ;
        RECT 28.000 20.720 30.520 21.280 ;
      LAYER met2 ;
        RECT 30.520 20.720 31.920 21.280 ;
      LAYER met2 ;
        RECT 31.920 21.000 41.720 21.280 ;
      LAYER met2 ;
        RECT 41.720 21.000 42.280 21.280 ;
      LAYER met2 ;
        RECT 31.920 20.720 41.440 21.000 ;
      LAYER met2 ;
        RECT 41.440 20.720 42.280 21.000 ;
      LAYER met2 ;
        RECT 42.280 20.720 43.960 21.280 ;
      LAYER met2 ;
        RECT 43.960 20.720 44.800 21.280 ;
      LAYER met2 ;
        RECT 44.800 21.000 45.360 21.560 ;
      LAYER met2 ;
        RECT 45.360 21.000 46.200 21.560 ;
      LAYER met2 ;
        RECT 46.200 21.000 46.480 21.560 ;
      LAYER met2 ;
        RECT 46.480 21.000 47.600 21.560 ;
      LAYER met2 ;
        RECT 47.600 21.280 48.720 21.560 ;
      LAYER met2 ;
        RECT 48.720 21.280 50.120 21.560 ;
      LAYER met2 ;
        RECT 47.600 21.000 48.440 21.280 ;
      LAYER met2 ;
        RECT 48.440 21.000 49.280 21.280 ;
      LAYER met2 ;
        RECT 49.280 21.000 49.560 21.280 ;
      LAYER met2 ;
        RECT 49.560 21.000 50.120 21.280 ;
      LAYER met2 ;
        RECT 50.120 21.000 50.680 21.560 ;
      LAYER met2 ;
        RECT 50.680 21.280 51.520 21.560 ;
      LAYER met2 ;
        RECT 51.520 21.280 52.080 21.560 ;
      LAYER met2 ;
        RECT 52.080 21.280 52.640 21.560 ;
      LAYER met2 ;
        RECT 52.640 21.280 55.720 21.560 ;
      LAYER met2 ;
        RECT 55.720 21.280 56.560 21.840 ;
      LAYER met2 ;
        RECT 56.560 21.560 70.840 21.840 ;
      LAYER met2 ;
        RECT 70.840 21.560 73.080 21.840 ;
      LAYER met2 ;
        RECT 73.080 21.560 79.520 21.840 ;
      LAYER met2 ;
        RECT 79.520 21.560 80.920 21.840 ;
      LAYER met2 ;
        RECT 80.920 21.560 90.160 21.840 ;
      LAYER met2 ;
        RECT 90.160 21.560 91.840 21.840 ;
      LAYER met2 ;
        RECT 56.560 21.280 70.000 21.560 ;
      LAYER met2 ;
        RECT 70.000 21.280 73.360 21.560 ;
      LAYER met2 ;
        RECT 73.360 21.280 77.560 21.560 ;
      LAYER met2 ;
        RECT 77.560 21.280 78.400 21.560 ;
      LAYER met2 ;
        RECT 78.400 21.280 79.520 21.560 ;
      LAYER met2 ;
        RECT 50.680 21.000 51.800 21.280 ;
      LAYER met2 ;
        RECT 51.800 21.000 52.360 21.280 ;
        RECT 44.800 20.720 45.080 21.000 ;
      LAYER met2 ;
        RECT 45.080 20.720 47.600 21.000 ;
      LAYER met2 ;
        RECT 47.600 20.720 48.160 21.000 ;
      LAYER met2 ;
        RECT 48.160 20.720 49.000 21.000 ;
      LAYER met2 ;
        RECT 49.000 20.720 49.560 21.000 ;
      LAYER met2 ;
        RECT 49.560 20.720 52.080 21.000 ;
      LAYER met2 ;
        RECT 52.080 20.720 52.360 21.000 ;
      LAYER met2 ;
        RECT 52.360 20.720 52.920 21.280 ;
      LAYER met2 ;
        RECT 52.920 21.000 56.000 21.280 ;
      LAYER met2 ;
        RECT 56.000 21.000 56.840 21.280 ;
      LAYER met2 ;
        RECT 56.840 21.000 68.880 21.280 ;
      LAYER met2 ;
        RECT 68.880 21.000 73.080 21.280 ;
      LAYER met2 ;
        RECT 73.080 21.000 77.560 21.280 ;
        RECT 52.920 20.720 56.280 21.000 ;
        RECT 0.000 20.160 4.760 20.720 ;
        RECT 0.000 19.600 0.840 20.160 ;
      LAYER met2 ;
        RECT 0.840 19.600 1.960 20.160 ;
      LAYER met2 ;
        RECT 0.000 17.640 0.560 19.600 ;
      LAYER met2 ;
        RECT 0.560 19.320 1.960 19.600 ;
      LAYER met2 ;
        RECT 1.960 19.320 4.760 20.160 ;
      LAYER met2 ;
        RECT 4.760 19.320 7.000 20.720 ;
      LAYER met2 ;
        RECT 7.000 20.440 13.160 20.720 ;
      LAYER met2 ;
        RECT 13.160 20.440 14.560 20.720 ;
      LAYER met2 ;
        RECT 7.000 19.320 13.440 20.440 ;
      LAYER met2 ;
        RECT 13.440 19.600 14.560 20.440 ;
      LAYER met2 ;
        RECT 14.560 20.160 18.480 20.720 ;
      LAYER met2 ;
        RECT 18.480 20.160 19.600 20.720 ;
      LAYER met2 ;
        RECT 19.600 20.440 22.680 20.720 ;
      LAYER met2 ;
        RECT 22.680 20.440 24.640 20.720 ;
      LAYER met2 ;
        RECT 24.640 20.440 26.320 20.720 ;
        RECT 14.560 19.600 18.200 20.160 ;
      LAYER met2 ;
        RECT 18.200 19.600 19.600 20.160 ;
      LAYER met2 ;
        RECT 19.600 19.600 22.400 20.440 ;
      LAYER met2 ;
        RECT 13.440 19.320 14.840 19.600 ;
        RECT 0.560 17.920 1.680 19.320 ;
      LAYER met2 ;
        RECT 1.680 17.920 4.760 19.320 ;
      LAYER met2 ;
        RECT 0.560 17.640 1.960 17.920 ;
      LAYER met2 ;
        RECT 0.000 16.240 0.840 17.640 ;
      LAYER met2 ;
        RECT 0.840 16.800 1.960 17.640 ;
      LAYER met2 ;
        RECT 1.960 16.800 4.760 17.920 ;
      LAYER met2 ;
        RECT 4.760 17.360 12.320 19.320 ;
      LAYER met2 ;
        RECT 12.320 17.640 13.720 19.320 ;
      LAYER met2 ;
        RECT 13.720 17.640 14.840 19.320 ;
      LAYER met2 ;
        RECT 12.320 17.360 13.440 17.640 ;
      LAYER met2 ;
        RECT 13.440 17.360 14.840 17.640 ;
      LAYER met2 ;
        RECT 14.840 17.360 18.200 19.600 ;
      LAYER met2 ;
        RECT 18.200 17.360 19.320 19.600 ;
      LAYER met2 ;
        RECT 19.320 19.040 22.400 19.600 ;
      LAYER met2 ;
        RECT 22.400 19.320 24.360 20.440 ;
      LAYER met2 ;
        RECT 24.360 19.320 26.320 20.440 ;
      LAYER met2 ;
        RECT 26.320 19.880 28.280 20.720 ;
      LAYER met2 ;
        RECT 28.280 19.880 30.800 20.720 ;
      LAYER met2 ;
        RECT 30.800 20.440 31.920 20.720 ;
      LAYER met2 ;
        RECT 31.920 20.440 41.160 20.720 ;
      LAYER met2 ;
        RECT 41.160 20.440 42.000 20.720 ;
      LAYER met2 ;
        RECT 42.000 20.440 43.680 20.720 ;
      LAYER met2 ;
        RECT 43.680 20.440 46.760 20.720 ;
      LAYER met2 ;
        RECT 46.760 20.440 47.040 20.720 ;
      LAYER met2 ;
        RECT 47.040 20.440 47.600 20.720 ;
      LAYER met2 ;
        RECT 47.600 20.440 47.880 20.720 ;
      LAYER met2 ;
        RECT 47.880 20.440 48.720 20.720 ;
      LAYER met2 ;
        RECT 48.720 20.440 49.560 20.720 ;
      LAYER met2 ;
        RECT 49.560 20.440 50.960 20.720 ;
      LAYER met2 ;
        RECT 50.960 20.440 51.520 20.720 ;
      LAYER met2 ;
        RECT 51.520 20.440 53.200 20.720 ;
      LAYER met2 ;
        RECT 53.200 20.440 54.040 20.720 ;
      LAYER met2 ;
        RECT 54.040 20.440 54.320 20.720 ;
      LAYER met2 ;
        RECT 54.320 20.440 56.280 20.720 ;
      LAYER met2 ;
        RECT 30.800 19.880 32.200 20.440 ;
      LAYER met2 ;
        RECT 32.200 20.160 41.160 20.440 ;
      LAYER met2 ;
        RECT 41.160 20.160 41.720 20.440 ;
      LAYER met2 ;
        RECT 41.720 20.160 43.400 20.440 ;
      LAYER met2 ;
        RECT 43.400 20.160 45.360 20.440 ;
      LAYER met2 ;
        RECT 45.360 20.160 45.640 20.440 ;
      LAYER met2 ;
        RECT 22.400 19.040 24.640 19.320 ;
      LAYER met2 ;
        RECT 24.640 19.040 26.320 19.320 ;
      LAYER met2 ;
        RECT 26.320 19.040 28.560 19.880 ;
      LAYER met2 ;
        RECT 19.320 18.480 22.680 19.040 ;
      LAYER met2 ;
        RECT 22.680 18.760 24.920 19.040 ;
      LAYER met2 ;
        RECT 24.920 18.760 26.040 19.040 ;
      LAYER met2 ;
        RECT 26.040 18.760 28.560 19.040 ;
        RECT 22.680 18.480 28.560 18.760 ;
      LAYER met2 ;
        RECT 19.320 17.920 22.960 18.480 ;
      LAYER met2 ;
        RECT 22.960 18.200 28.560 18.480 ;
      LAYER met2 ;
        RECT 28.560 18.200 31.080 19.880 ;
      LAYER met2 ;
        RECT 22.960 17.920 28.280 18.200 ;
      LAYER met2 ;
        RECT 19.320 17.640 23.240 17.920 ;
      LAYER met2 ;
        RECT 23.240 17.640 28.280 17.920 ;
      LAYER met2 ;
        RECT 19.320 17.360 23.800 17.640 ;
      LAYER met2 ;
        RECT 23.800 17.360 25.760 17.640 ;
      LAYER met2 ;
        RECT 25.760 17.360 26.320 17.640 ;
      LAYER met2 ;
        RECT 26.320 17.360 28.280 17.640 ;
      LAYER met2 ;
        RECT 28.280 17.360 31.080 18.200 ;
      LAYER met2 ;
        RECT 31.080 17.360 32.200 19.880 ;
      LAYER met2 ;
        RECT 32.200 19.040 40.880 20.160 ;
      LAYER met2 ;
        RECT 40.880 19.880 41.720 20.160 ;
      LAYER met2 ;
        RECT 41.720 19.880 43.120 20.160 ;
      LAYER met2 ;
        RECT 43.120 19.880 45.080 20.160 ;
      LAYER met2 ;
        RECT 45.080 19.880 45.640 20.160 ;
      LAYER met2 ;
        RECT 45.640 19.880 46.480 20.440 ;
      LAYER met2 ;
        RECT 46.480 19.880 47.040 20.440 ;
      LAYER met2 ;
        RECT 47.040 20.160 48.440 20.440 ;
      LAYER met2 ;
        RECT 48.440 20.160 49.560 20.440 ;
      LAYER met2 ;
        RECT 49.560 20.160 50.400 20.440 ;
      LAYER met2 ;
        RECT 50.400 20.160 52.080 20.440 ;
      LAYER met2 ;
        RECT 52.080 20.160 53.480 20.440 ;
      LAYER met2 ;
        RECT 53.480 20.160 54.040 20.440 ;
      LAYER met2 ;
        RECT 54.040 20.160 54.600 20.440 ;
      LAYER met2 ;
        RECT 54.600 20.160 56.280 20.440 ;
      LAYER met2 ;
        RECT 56.280 20.160 56.840 21.000 ;
      LAYER met2 ;
        RECT 56.840 20.160 67.760 21.000 ;
      LAYER met2 ;
        RECT 67.760 20.720 72.800 21.000 ;
      LAYER met2 ;
        RECT 72.800 20.720 77.560 21.000 ;
      LAYER met2 ;
        RECT 47.040 19.880 48.160 20.160 ;
      LAYER met2 ;
        RECT 48.160 19.880 52.360 20.160 ;
      LAYER met2 ;
        RECT 52.360 19.880 53.480 20.160 ;
      LAYER met2 ;
        RECT 53.480 19.880 54.320 20.160 ;
      LAYER met2 ;
        RECT 54.320 19.880 54.600 20.160 ;
      LAYER met2 ;
        RECT 54.600 19.880 56.560 20.160 ;
      LAYER met2 ;
        RECT 40.880 19.320 41.440 19.880 ;
      LAYER met2 ;
        RECT 41.440 19.600 42.840 19.880 ;
      LAYER met2 ;
        RECT 42.840 19.600 44.800 19.880 ;
      LAYER met2 ;
        RECT 44.800 19.600 45.640 19.880 ;
      LAYER met2 ;
        RECT 45.640 19.600 46.200 19.880 ;
      LAYER met2 ;
        RECT 46.200 19.600 47.320 19.880 ;
        RECT 41.440 19.320 41.720 19.600 ;
      LAYER met2 ;
        RECT 41.720 19.320 42.280 19.600 ;
      LAYER met2 ;
        RECT 42.280 19.320 42.560 19.600 ;
      LAYER met2 ;
        RECT 42.560 19.320 43.680 19.600 ;
        RECT 40.880 19.040 43.680 19.320 ;
      LAYER met2 ;
        RECT 32.200 18.480 41.160 19.040 ;
      LAYER met2 ;
        RECT 41.160 18.760 42.560 19.040 ;
        RECT 41.160 18.480 41.720 18.760 ;
      LAYER met2 ;
        RECT 41.720 18.480 42.000 18.760 ;
        RECT 32.200 18.200 42.000 18.480 ;
      LAYER met2 ;
        RECT 42.000 18.200 42.560 18.760 ;
      LAYER met2 ;
        RECT 42.560 18.200 42.840 19.040 ;
        RECT 32.200 17.360 41.720 18.200 ;
      LAYER met2 ;
        RECT 41.720 17.360 42.280 18.200 ;
      LAYER met2 ;
        RECT 42.280 17.360 42.840 18.200 ;
      LAYER met2 ;
        RECT 42.840 17.920 43.680 19.040 ;
      LAYER met2 ;
        RECT 43.680 17.920 43.960 19.600 ;
      LAYER met2 ;
        RECT 42.840 17.360 43.400 17.920 ;
        RECT 0.840 16.240 2.240 16.800 ;
      LAYER met2 ;
        RECT 0.000 15.680 1.120 16.240 ;
      LAYER met2 ;
        RECT 1.120 15.960 2.240 16.240 ;
      LAYER met2 ;
        RECT 2.240 15.960 4.760 16.800 ;
      LAYER met2 ;
        RECT 4.760 15.960 7.000 17.360 ;
      LAYER met2 ;
        RECT 7.000 15.960 8.120 17.360 ;
      LAYER met2 ;
        RECT 1.120 15.680 2.520 15.960 ;
      LAYER met2 ;
        RECT 2.520 15.680 8.120 15.960 ;
        RECT 0.000 15.120 1.400 15.680 ;
      LAYER met2 ;
        RECT 1.400 15.120 2.800 15.680 ;
      LAYER met2 ;
        RECT 2.800 15.120 8.120 15.680 ;
        RECT 0.000 14.560 1.680 15.120 ;
      LAYER met2 ;
        RECT 1.680 14.840 3.080 15.120 ;
      LAYER met2 ;
        RECT 3.080 14.840 8.120 15.120 ;
      LAYER met2 ;
        RECT 1.680 14.560 3.360 14.840 ;
      LAYER met2 ;
        RECT 3.360 14.560 8.120 14.840 ;
        RECT 0.000 14.280 1.960 14.560 ;
      LAYER met2 ;
        RECT 1.960 14.280 3.640 14.560 ;
      LAYER met2 ;
        RECT 3.640 14.280 8.120 14.560 ;
        RECT 0.000 14.000 2.240 14.280 ;
      LAYER met2 ;
        RECT 2.240 14.000 3.920 14.280 ;
      LAYER met2 ;
        RECT 3.920 14.000 8.120 14.280 ;
        RECT 0.000 13.720 2.520 14.000 ;
      LAYER met2 ;
        RECT 2.520 13.720 4.200 14.000 ;
      LAYER met2 ;
        RECT 4.200 13.720 8.120 14.000 ;
        RECT 0.000 13.440 2.800 13.720 ;
      LAYER met2 ;
        RECT 2.800 13.440 4.480 13.720 ;
      LAYER met2 ;
        RECT 4.480 13.440 8.120 13.720 ;
        RECT 0.000 13.160 3.080 13.440 ;
      LAYER met2 ;
        RECT 3.080 13.160 5.040 13.440 ;
      LAYER met2 ;
        RECT 5.040 13.160 8.120 13.440 ;
        RECT 0.000 12.880 3.360 13.160 ;
      LAYER met2 ;
        RECT 3.360 12.880 5.600 13.160 ;
      LAYER met2 ;
        RECT 5.600 12.880 8.120 13.160 ;
        RECT 0.000 12.600 3.640 12.880 ;
      LAYER met2 ;
        RECT 3.640 12.600 7.000 12.880 ;
      LAYER met2 ;
        RECT 7.000 12.600 8.120 12.880 ;
      LAYER met2 ;
        RECT 8.120 12.600 10.360 17.360 ;
      LAYER met2 ;
        RECT 10.360 16.800 13.440 17.360 ;
      LAYER met2 ;
        RECT 13.440 16.800 14.560 17.360 ;
      LAYER met2 ;
        RECT 14.560 16.800 18.200 17.360 ;
      LAYER met2 ;
        RECT 18.200 16.800 19.600 17.360 ;
      LAYER met2 ;
        RECT 19.600 17.080 26.320 17.360 ;
      LAYER met2 ;
        RECT 26.320 17.080 28.000 17.360 ;
      LAYER met2 ;
        RECT 19.600 16.800 26.040 17.080 ;
      LAYER met2 ;
        RECT 26.040 16.800 28.000 17.080 ;
      LAYER met2 ;
        RECT 28.000 16.800 30.800 17.360 ;
      LAYER met2 ;
        RECT 30.800 16.800 32.200 17.360 ;
      LAYER met2 ;
        RECT 32.200 16.800 41.440 17.360 ;
      LAYER met2 ;
        RECT 41.440 17.080 42.280 17.360 ;
      LAYER met2 ;
        RECT 42.280 17.080 42.560 17.360 ;
      LAYER met2 ;
        RECT 42.560 17.080 43.400 17.360 ;
      LAYER met2 ;
        RECT 43.400 17.080 43.960 17.920 ;
        RECT 10.360 15.960 13.160 16.800 ;
      LAYER met2 ;
        RECT 13.160 16.240 14.560 16.800 ;
      LAYER met2 ;
        RECT 14.560 16.240 18.480 16.800 ;
      LAYER met2 ;
        RECT 18.480 16.520 19.600 16.800 ;
      LAYER met2 ;
        RECT 19.600 16.520 25.760 16.800 ;
      LAYER met2 ;
        RECT 25.760 16.520 27.720 16.800 ;
        RECT 13.160 15.960 14.280 16.240 ;
      LAYER met2 ;
        RECT 14.280 15.960 18.480 16.240 ;
      LAYER met2 ;
        RECT 18.480 15.960 19.880 16.520 ;
      LAYER met2 ;
        RECT 19.880 16.240 25.200 16.520 ;
      LAYER met2 ;
        RECT 25.200 16.240 27.720 16.520 ;
      LAYER met2 ;
        RECT 27.720 16.240 30.800 16.800 ;
      LAYER met2 ;
        RECT 30.800 16.240 31.920 16.800 ;
      LAYER met2 ;
        RECT 19.880 15.960 24.360 16.240 ;
      LAYER met2 ;
        RECT 24.360 15.960 27.440 16.240 ;
      LAYER met2 ;
        RECT 27.440 15.960 30.520 16.240 ;
      LAYER met2 ;
        RECT 30.520 15.960 31.920 16.240 ;
      LAYER met2 ;
        RECT 31.920 15.960 41.440 16.800 ;
      LAYER met2 ;
        RECT 41.440 15.960 42.000 17.080 ;
      LAYER met2 ;
        RECT 42.000 16.800 42.560 17.080 ;
      LAYER met2 ;
        RECT 42.560 16.800 43.120 17.080 ;
      LAYER met2 ;
        RECT 42.000 15.960 42.280 16.800 ;
      LAYER met2 ;
        RECT 42.280 16.240 43.120 16.800 ;
      LAYER met2 ;
        RECT 43.120 16.240 43.960 17.080 ;
      LAYER met2 ;
        RECT 42.280 15.960 42.840 16.240 ;
      LAYER met2 ;
        RECT 10.360 15.400 12.880 15.960 ;
      LAYER met2 ;
        RECT 12.880 15.680 14.280 15.960 ;
      LAYER met2 ;
        RECT 14.280 15.680 18.760 15.960 ;
      LAYER met2 ;
        RECT 18.760 15.680 19.880 15.960 ;
      LAYER met2 ;
        RECT 19.880 15.680 23.240 15.960 ;
      LAYER met2 ;
        RECT 23.240 15.680 27.160 15.960 ;
      LAYER met2 ;
        RECT 27.160 15.680 30.520 15.960 ;
      LAYER met2 ;
        RECT 30.520 15.680 31.640 15.960 ;
        RECT 12.880 15.400 14.000 15.680 ;
      LAYER met2 ;
        RECT 14.000 15.400 18.760 15.680 ;
      LAYER met2 ;
        RECT 18.760 15.400 20.160 15.680 ;
      LAYER met2 ;
        RECT 20.160 15.400 23.240 15.680 ;
      LAYER met2 ;
        RECT 23.240 15.400 26.880 15.680 ;
      LAYER met2 ;
        RECT 26.880 15.400 30.240 15.680 ;
      LAYER met2 ;
        RECT 30.240 15.400 31.640 15.680 ;
      LAYER met2 ;
        RECT 31.640 15.400 41.440 15.960 ;
      LAYER met2 ;
        RECT 41.440 15.400 42.840 15.960 ;
      LAYER met2 ;
        RECT 42.840 15.400 43.960 16.240 ;
      LAYER met2 ;
        RECT 43.960 15.400 44.520 19.600 ;
      LAYER met2 ;
        RECT 44.520 19.320 47.320 19.600 ;
      LAYER met2 ;
        RECT 47.320 19.320 48.160 19.880 ;
      LAYER met2 ;
        RECT 48.160 19.600 52.640 19.880 ;
      LAYER met2 ;
        RECT 52.640 19.600 53.760 19.880 ;
      LAYER met2 ;
        RECT 53.760 19.600 54.320 19.880 ;
      LAYER met2 ;
        RECT 54.320 19.600 54.880 19.880 ;
      LAYER met2 ;
        RECT 48.160 19.320 52.920 19.600 ;
      LAYER met2 ;
        RECT 52.920 19.320 54.040 19.600 ;
      LAYER met2 ;
        RECT 54.040 19.320 54.600 19.600 ;
        RECT 44.520 18.760 47.600 19.320 ;
      LAYER met2 ;
        RECT 47.600 18.760 47.880 19.320 ;
      LAYER met2 ;
        RECT 47.880 18.760 50.960 19.320 ;
      LAYER met2 ;
        RECT 50.960 19.040 51.240 19.320 ;
      LAYER met2 ;
        RECT 51.240 19.040 52.920 19.320 ;
      LAYER met2 ;
        RECT 52.920 19.040 54.320 19.320 ;
      LAYER met2 ;
        RECT 54.320 19.040 54.600 19.320 ;
      LAYER met2 ;
        RECT 54.600 19.040 54.880 19.600 ;
      LAYER met2 ;
        RECT 10.360 15.120 12.600 15.400 ;
      LAYER met2 ;
        RECT 12.600 15.120 14.000 15.400 ;
      LAYER met2 ;
        RECT 14.000 15.120 19.040 15.400 ;
        RECT 10.360 14.840 12.320 15.120 ;
      LAYER met2 ;
        RECT 12.320 14.840 13.720 15.120 ;
      LAYER met2 ;
        RECT 13.720 14.840 19.040 15.120 ;
      LAYER met2 ;
        RECT 19.040 14.840 20.440 15.400 ;
      LAYER met2 ;
        RECT 20.440 14.840 23.240 15.400 ;
      LAYER met2 ;
        RECT 23.240 15.120 26.600 15.400 ;
      LAYER met2 ;
        RECT 26.600 15.120 29.960 15.400 ;
      LAYER met2 ;
        RECT 23.240 14.840 26.040 15.120 ;
      LAYER met2 ;
        RECT 26.040 14.840 29.960 15.120 ;
      LAYER met2 ;
        RECT 29.960 14.840 31.360 15.400 ;
      LAYER met2 ;
        RECT 31.360 15.120 41.440 15.400 ;
      LAYER met2 ;
        RECT 41.440 15.120 43.120 15.400 ;
      LAYER met2 ;
        RECT 43.120 15.120 44.240 15.400 ;
      LAYER met2 ;
        RECT 44.240 15.120 44.520 15.400 ;
      LAYER met2 ;
        RECT 44.520 15.120 50.960 18.760 ;
      LAYER met2 ;
        RECT 50.960 15.120 51.520 19.040 ;
      LAYER met2 ;
        RECT 51.520 18.480 52.920 19.040 ;
      LAYER met2 ;
        RECT 52.920 18.760 54.880 19.040 ;
        RECT 52.920 18.480 53.760 18.760 ;
      LAYER met2 ;
        RECT 53.760 18.480 54.040 18.760 ;
      LAYER met2 ;
        RECT 54.040 18.480 54.880 18.760 ;
      LAYER met2 ;
        RECT 51.520 17.080 53.200 18.480 ;
      LAYER met2 ;
        RECT 53.200 17.080 53.760 18.480 ;
      LAYER met2 ;
        RECT 53.760 17.920 54.320 18.480 ;
      LAYER met2 ;
        RECT 54.320 17.920 54.880 18.480 ;
      LAYER met2 ;
        RECT 54.880 17.920 56.560 19.880 ;
      LAYER met2 ;
        RECT 56.560 18.200 57.120 20.160 ;
      LAYER met2 ;
        RECT 57.120 19.600 67.760 20.160 ;
      LAYER met2 ;
        RECT 67.760 19.880 72.240 20.720 ;
        RECT 67.760 19.600 69.720 19.880 ;
      LAYER met2 ;
        RECT 69.720 19.600 70.560 19.880 ;
        RECT 57.120 19.040 70.560 19.600 ;
      LAYER met2 ;
        RECT 70.560 19.320 72.240 19.880 ;
      LAYER met2 ;
        RECT 72.240 19.320 77.560 20.720 ;
      LAYER met2 ;
        RECT 70.560 19.040 74.200 19.320 ;
      LAYER met2 ;
        RECT 57.120 18.200 67.200 19.040 ;
      LAYER met2 ;
        RECT 56.560 17.920 57.400 18.200 ;
      LAYER met2 ;
        RECT 53.760 17.360 56.840 17.920 ;
      LAYER met2 ;
        RECT 56.840 17.360 57.400 17.920 ;
      LAYER met2 ;
        RECT 57.400 17.640 67.200 18.200 ;
      LAYER met2 ;
        RECT 67.200 17.640 74.200 19.040 ;
      LAYER met2 ;
        RECT 74.200 18.760 77.560 19.320 ;
      LAYER met2 ;
        RECT 77.560 18.760 79.240 21.280 ;
      LAYER met2 ;
        RECT 74.200 17.920 77.280 18.760 ;
      LAYER met2 ;
        RECT 77.280 18.200 79.240 18.760 ;
      LAYER met2 ;
        RECT 79.240 18.200 79.520 21.280 ;
      LAYER met2 ;
        RECT 77.280 17.920 78.960 18.200 ;
      LAYER met2 ;
        RECT 74.200 17.640 77.000 17.920 ;
        RECT 57.400 17.360 70.280 17.640 ;
        RECT 53.760 17.080 57.120 17.360 ;
        RECT 51.520 15.960 52.920 17.080 ;
      LAYER met2 ;
        RECT 52.920 15.960 53.480 17.080 ;
      LAYER met2 ;
        RECT 53.480 16.800 57.120 17.080 ;
      LAYER met2 ;
        RECT 57.120 16.800 57.680 17.360 ;
      LAYER met2 ;
        RECT 57.680 16.800 70.280 17.360 ;
      LAYER met2 ;
        RECT 70.280 17.080 72.240 17.640 ;
      LAYER met2 ;
        RECT 72.240 17.360 77.000 17.640 ;
      LAYER met2 ;
        RECT 77.000 17.360 78.960 17.920 ;
      LAYER met2 ;
        RECT 72.240 17.080 76.720 17.360 ;
      LAYER met2 ;
        RECT 76.720 17.080 78.960 17.360 ;
      LAYER met2 ;
        RECT 78.960 17.080 79.520 18.200 ;
      LAYER met2 ;
        RECT 79.520 17.080 81.200 21.560 ;
      LAYER met2 ;
        RECT 81.200 19.880 89.880 21.560 ;
      LAYER met2 ;
        RECT 89.880 19.880 91.840 21.560 ;
      LAYER met2 ;
        RECT 91.840 19.880 92.400 21.840 ;
        RECT 81.200 19.040 89.600 19.880 ;
      LAYER met2 ;
        RECT 89.600 19.040 91.560 19.880 ;
      LAYER met2 ;
        RECT 91.560 19.040 92.400 19.880 ;
        RECT 81.200 18.760 89.320 19.040 ;
        RECT 81.200 18.480 82.880 18.760 ;
      LAYER met2 ;
        RECT 82.880 18.480 83.440 18.760 ;
      LAYER met2 ;
        RECT 83.440 18.480 89.320 18.760 ;
      LAYER met2 ;
        RECT 89.320 18.480 91.280 19.040 ;
      LAYER met2 ;
        RECT 81.200 17.920 82.600 18.480 ;
      LAYER met2 ;
        RECT 82.600 18.200 83.720 18.480 ;
      LAYER met2 ;
        RECT 83.720 18.200 89.040 18.480 ;
      LAYER met2 ;
        RECT 89.040 18.200 91.280 18.480 ;
      LAYER met2 ;
        RECT 91.280 18.200 92.400 19.040 ;
      LAYER met2 ;
        RECT 82.600 17.920 84.280 18.200 ;
      LAYER met2 ;
        RECT 84.280 17.920 88.760 18.200 ;
      LAYER met2 ;
        RECT 88.760 17.920 91.000 18.200 ;
      LAYER met2 ;
        RECT 81.200 17.640 82.320 17.920 ;
      LAYER met2 ;
        RECT 82.320 17.640 84.560 17.920 ;
      LAYER met2 ;
        RECT 84.560 17.640 88.480 17.920 ;
      LAYER met2 ;
        RECT 88.480 17.640 91.000 17.920 ;
      LAYER met2 ;
        RECT 91.000 17.640 92.400 18.200 ;
        RECT 81.200 17.360 82.040 17.640 ;
      LAYER met2 ;
        RECT 82.040 17.360 84.560 17.640 ;
      LAYER met2 ;
        RECT 84.560 17.360 88.200 17.640 ;
      LAYER met2 ;
        RECT 88.200 17.360 90.720 17.640 ;
      LAYER met2 ;
        RECT 90.720 17.360 92.400 17.640 ;
        RECT 81.200 17.080 81.760 17.360 ;
      LAYER met2 ;
        RECT 81.760 17.080 84.280 17.360 ;
      LAYER met2 ;
        RECT 84.280 17.080 87.920 17.360 ;
      LAYER met2 ;
        RECT 87.920 17.080 90.440 17.360 ;
        RECT 70.280 16.800 71.960 17.080 ;
      LAYER met2 ;
        RECT 53.480 16.240 57.400 16.800 ;
      LAYER met2 ;
        RECT 57.400 16.240 57.960 16.800 ;
      LAYER met2 ;
        RECT 57.960 16.520 70.000 16.800 ;
      LAYER met2 ;
        RECT 70.000 16.520 71.960 16.800 ;
      LAYER met2 ;
        RECT 71.960 16.520 76.440 17.080 ;
      LAYER met2 ;
        RECT 76.440 16.800 78.680 17.080 ;
      LAYER met2 ;
        RECT 78.680 16.800 79.520 17.080 ;
      LAYER met2 ;
        RECT 79.520 16.800 84.000 17.080 ;
      LAYER met2 ;
        RECT 84.000 16.800 87.640 17.080 ;
      LAYER met2 ;
        RECT 87.640 16.800 90.440 17.080 ;
      LAYER met2 ;
        RECT 90.440 16.800 92.400 17.360 ;
      LAYER met2 ;
        RECT 76.440 16.520 78.400 16.800 ;
      LAYER met2 ;
        RECT 57.960 16.240 69.720 16.520 ;
      LAYER met2 ;
        RECT 69.720 16.240 71.680 16.520 ;
      LAYER met2 ;
        RECT 71.680 16.240 76.160 16.520 ;
      LAYER met2 ;
        RECT 76.160 16.240 78.400 16.520 ;
      LAYER met2 ;
        RECT 78.400 16.240 79.520 16.800 ;
      LAYER met2 ;
        RECT 79.520 16.520 83.720 16.800 ;
      LAYER met2 ;
        RECT 83.720 16.520 87.360 16.800 ;
      LAYER met2 ;
        RECT 87.360 16.520 90.160 16.800 ;
      LAYER met2 ;
        RECT 90.160 16.520 92.400 16.800 ;
      LAYER met2 ;
        RECT 79.520 16.240 83.440 16.520 ;
      LAYER met2 ;
        RECT 83.440 16.240 86.800 16.520 ;
      LAYER met2 ;
        RECT 86.800 16.240 89.880 16.520 ;
      LAYER met2 ;
        RECT 89.880 16.240 92.400 16.520 ;
        RECT 53.480 15.960 57.680 16.240 ;
        RECT 51.520 15.120 52.640 15.960 ;
        RECT 31.360 14.840 41.160 15.120 ;
      LAYER met2 ;
        RECT 41.160 14.840 42.000 15.120 ;
      LAYER met2 ;
        RECT 42.000 14.840 42.560 15.120 ;
      LAYER met2 ;
        RECT 42.560 14.840 43.400 15.120 ;
      LAYER met2 ;
        RECT 43.400 14.840 52.640 15.120 ;
        RECT 10.360 14.560 12.040 14.840 ;
      LAYER met2 ;
        RECT 12.040 14.560 13.720 14.840 ;
      LAYER met2 ;
        RECT 13.720 14.560 19.320 14.840 ;
      LAYER met2 ;
        RECT 19.320 14.560 20.720 14.840 ;
      LAYER met2 ;
        RECT 20.720 14.560 23.240 14.840 ;
      LAYER met2 ;
        RECT 23.240 14.560 25.480 14.840 ;
      LAYER met2 ;
        RECT 25.480 14.560 29.680 14.840 ;
      LAYER met2 ;
        RECT 29.680 14.560 31.080 14.840 ;
      LAYER met2 ;
        RECT 31.080 14.560 41.160 14.840 ;
      LAYER met2 ;
        RECT 41.160 14.560 41.720 14.840 ;
      LAYER met2 ;
        RECT 10.360 14.280 11.760 14.560 ;
      LAYER met2 ;
        RECT 11.760 14.280 13.440 14.560 ;
      LAYER met2 ;
        RECT 13.440 14.280 19.600 14.560 ;
      LAYER met2 ;
        RECT 19.600 14.280 21.000 14.560 ;
      LAYER met2 ;
        RECT 21.000 14.280 29.400 14.560 ;
      LAYER met2 ;
        RECT 29.400 14.280 31.080 14.560 ;
      LAYER met2 ;
        RECT 31.080 14.280 40.880 14.560 ;
      LAYER met2 ;
        RECT 40.880 14.280 41.720 14.560 ;
      LAYER met2 ;
        RECT 41.720 14.280 42.560 14.840 ;
      LAYER met2 ;
        RECT 42.560 14.560 43.680 14.840 ;
      LAYER met2 ;
        RECT 43.680 14.560 52.640 14.840 ;
      LAYER met2 ;
        RECT 52.640 14.560 53.200 15.960 ;
      LAYER met2 ;
        RECT 53.200 15.680 57.680 15.960 ;
        RECT 53.200 14.560 55.440 15.680 ;
      LAYER met2 ;
        RECT 55.440 15.120 55.720 15.680 ;
      LAYER met2 ;
        RECT 55.720 15.400 57.680 15.680 ;
        RECT 55.720 15.120 56.840 15.400 ;
      LAYER met2 ;
        RECT 56.840 15.120 57.120 15.400 ;
      LAYER met2 ;
        RECT 57.120 15.120 57.680 15.400 ;
      LAYER met2 ;
        RECT 42.560 14.280 43.960 14.560 ;
      LAYER met2 ;
        RECT 43.960 14.280 46.200 14.560 ;
        RECT 10.360 14.000 11.480 14.280 ;
      LAYER met2 ;
        RECT 11.480 14.000 13.160 14.280 ;
      LAYER met2 ;
        RECT 13.160 14.000 19.600 14.280 ;
      LAYER met2 ;
        RECT 19.600 14.000 21.280 14.280 ;
      LAYER met2 ;
        RECT 21.280 14.000 29.120 14.280 ;
      LAYER met2 ;
        RECT 29.120 14.000 30.800 14.280 ;
      LAYER met2 ;
        RECT 30.800 14.000 40.880 14.280 ;
        RECT 10.360 13.720 11.200 14.000 ;
      LAYER met2 ;
        RECT 11.200 13.720 12.880 14.000 ;
      LAYER met2 ;
        RECT 12.880 13.720 19.880 14.000 ;
      LAYER met2 ;
        RECT 19.880 13.720 21.560 14.000 ;
      LAYER met2 ;
        RECT 21.560 13.720 28.840 14.000 ;
      LAYER met2 ;
        RECT 28.840 13.720 30.520 14.000 ;
      LAYER met2 ;
        RECT 30.520 13.720 40.880 14.000 ;
      LAYER met2 ;
        RECT 40.880 13.720 42.280 14.280 ;
      LAYER met2 ;
        RECT 42.280 13.720 42.560 14.280 ;
      LAYER met2 ;
        RECT 42.560 13.720 43.120 14.280 ;
      LAYER met2 ;
        RECT 43.120 14.000 43.400 14.280 ;
      LAYER met2 ;
        RECT 43.400 14.000 44.520 14.280 ;
      LAYER met2 ;
        RECT 44.520 14.000 46.200 14.280 ;
      LAYER met2 ;
        RECT 46.200 14.000 50.400 14.560 ;
      LAYER met2 ;
        RECT 50.400 14.280 52.640 14.560 ;
      LAYER met2 ;
        RECT 52.640 14.280 53.480 14.560 ;
      LAYER met2 ;
        RECT 43.120 13.720 43.680 14.000 ;
      LAYER met2 ;
        RECT 43.680 13.720 44.800 14.000 ;
      LAYER met2 ;
        RECT 44.800 13.720 46.200 14.000 ;
      LAYER met2 ;
        RECT 46.200 13.720 46.760 14.000 ;
      LAYER met2 ;
        RECT 46.760 13.720 49.840 14.000 ;
        RECT 0.000 12.320 4.200 12.600 ;
      LAYER met2 ;
        RECT 4.200 12.320 10.360 12.600 ;
      LAYER met2 ;
        RECT 10.360 12.320 10.920 13.720 ;
      LAYER met2 ;
        RECT 10.920 13.440 12.600 13.720 ;
      LAYER met2 ;
        RECT 12.600 13.440 20.160 13.720 ;
      LAYER met2 ;
        RECT 20.160 13.440 22.120 13.720 ;
      LAYER met2 ;
        RECT 22.120 13.440 28.280 13.720 ;
      LAYER met2 ;
        RECT 28.280 13.440 30.240 13.720 ;
      LAYER met2 ;
        RECT 30.240 13.440 41.160 13.720 ;
      LAYER met2 ;
        RECT 41.160 13.440 43.120 13.720 ;
      LAYER met2 ;
        RECT 43.120 13.440 43.400 13.720 ;
      LAYER met2 ;
        RECT 43.400 13.440 45.640 13.720 ;
      LAYER met2 ;
        RECT 45.640 13.440 46.480 13.720 ;
      LAYER met2 ;
        RECT 10.920 13.160 12.320 13.440 ;
      LAYER met2 ;
        RECT 12.320 13.160 20.440 13.440 ;
      LAYER met2 ;
        RECT 20.440 13.160 22.680 13.440 ;
      LAYER met2 ;
        RECT 22.680 13.160 27.720 13.440 ;
      LAYER met2 ;
        RECT 27.720 13.160 29.960 13.440 ;
      LAYER met2 ;
        RECT 29.960 13.160 41.440 13.440 ;
      LAYER met2 ;
        RECT 41.440 13.160 46.200 13.440 ;
      LAYER met2 ;
        RECT 46.200 13.160 46.480 13.440 ;
      LAYER met2 ;
        RECT 46.480 13.160 47.040 13.720 ;
      LAYER met2 ;
        RECT 47.040 13.160 49.840 13.720 ;
      LAYER met2 ;
        RECT 10.920 12.880 12.040 13.160 ;
      LAYER met2 ;
        RECT 12.040 12.880 20.720 13.160 ;
      LAYER met2 ;
        RECT 20.720 12.880 23.240 13.160 ;
      LAYER met2 ;
        RECT 23.240 12.880 27.160 13.160 ;
      LAYER met2 ;
        RECT 27.160 12.880 29.680 13.160 ;
      LAYER met2 ;
        RECT 29.680 12.880 41.440 13.160 ;
      LAYER met2 ;
        RECT 41.440 12.880 47.320 13.160 ;
      LAYER met2 ;
        RECT 47.320 12.880 49.840 13.160 ;
      LAYER met2 ;
        RECT 49.840 12.880 50.400 14.000 ;
      LAYER met2 ;
        RECT 50.400 13.720 52.920 14.280 ;
      LAYER met2 ;
        RECT 52.920 13.720 53.480 14.280 ;
      LAYER met2 ;
        RECT 50.400 13.440 52.640 13.720 ;
      LAYER met2 ;
        RECT 52.640 13.440 53.480 13.720 ;
      LAYER met2 ;
        RECT 50.400 13.160 52.360 13.440 ;
      LAYER met2 ;
        RECT 52.360 13.160 53.480 13.440 ;
      LAYER met2 ;
        RECT 53.480 13.160 53.760 14.560 ;
      LAYER met2 ;
        RECT 53.760 14.280 54.320 14.560 ;
      LAYER met2 ;
        RECT 54.320 14.280 55.440 14.560 ;
      LAYER met2 ;
        RECT 53.760 13.160 54.880 14.280 ;
      LAYER met2 ;
        RECT 54.880 13.440 55.440 14.280 ;
      LAYER met2 ;
        RECT 55.440 13.720 56.000 15.120 ;
      LAYER met2 ;
        RECT 56.000 14.560 56.840 15.120 ;
      LAYER met2 ;
        RECT 56.840 14.840 57.400 15.120 ;
      LAYER met2 ;
        RECT 57.400 14.840 57.680 15.120 ;
      LAYER met2 ;
        RECT 57.680 14.840 58.240 16.240 ;
      LAYER met2 ;
        RECT 58.240 15.960 69.440 16.240 ;
      LAYER met2 ;
        RECT 69.440 15.960 71.680 16.240 ;
      LAYER met2 ;
        RECT 71.680 15.960 75.880 16.240 ;
        RECT 58.240 15.120 68.880 15.960 ;
      LAYER met2 ;
        RECT 68.880 15.680 71.400 15.960 ;
      LAYER met2 ;
        RECT 71.400 15.680 75.880 15.960 ;
      LAYER met2 ;
        RECT 75.880 15.680 78.120 16.240 ;
      LAYER met2 ;
        RECT 78.120 15.680 79.520 16.240 ;
      LAYER met2 ;
        RECT 79.520 15.960 83.160 16.240 ;
      LAYER met2 ;
        RECT 83.160 15.960 86.240 16.240 ;
      LAYER met2 ;
        RECT 86.240 15.960 89.600 16.240 ;
      LAYER met2 ;
        RECT 89.600 15.960 92.400 16.240 ;
      LAYER met2 ;
        RECT 79.520 15.680 82.880 15.960 ;
      LAYER met2 ;
        RECT 82.880 15.680 85.680 15.960 ;
      LAYER met2 ;
        RECT 85.680 15.680 89.320 15.960 ;
      LAYER met2 ;
        RECT 89.320 15.680 92.400 15.960 ;
      LAYER met2 ;
        RECT 68.880 15.400 71.120 15.680 ;
      LAYER met2 ;
        RECT 71.120 15.400 76.160 15.680 ;
      LAYER met2 ;
        RECT 76.160 15.400 77.840 15.680 ;
      LAYER met2 ;
        RECT 77.840 15.400 79.520 15.680 ;
      LAYER met2 ;
        RECT 79.520 15.400 82.320 15.680 ;
      LAYER met2 ;
        RECT 82.320 15.400 85.680 15.680 ;
      LAYER met2 ;
        RECT 85.680 15.400 88.760 15.680 ;
      LAYER met2 ;
        RECT 88.760 15.400 92.400 15.680 ;
      LAYER met2 ;
        RECT 68.880 15.120 70.840 15.400 ;
      LAYER met2 ;
        RECT 70.840 15.120 76.440 15.400 ;
      LAYER met2 ;
        RECT 76.440 15.120 77.560 15.400 ;
      LAYER met2 ;
        RECT 77.560 15.120 79.520 15.400 ;
      LAYER met2 ;
        RECT 79.520 15.120 81.760 15.400 ;
      LAYER met2 ;
        RECT 81.760 15.120 85.960 15.400 ;
      LAYER met2 ;
        RECT 85.960 15.120 88.200 15.400 ;
      LAYER met2 ;
        RECT 88.200 15.120 92.400 15.400 ;
        RECT 58.240 14.840 69.160 15.120 ;
      LAYER met2 ;
        RECT 69.160 14.840 70.560 15.120 ;
      LAYER met2 ;
        RECT 70.560 14.840 76.440 15.120 ;
      LAYER met2 ;
        RECT 76.440 14.840 77.000 15.120 ;
      LAYER met2 ;
        RECT 77.000 14.840 80.080 15.120 ;
      LAYER met2 ;
        RECT 80.080 14.840 80.920 15.120 ;
      LAYER met2 ;
        RECT 80.920 14.840 86.240 15.120 ;
      LAYER met2 ;
        RECT 86.240 14.840 87.640 15.120 ;
      LAYER met2 ;
        RECT 87.640 14.840 92.400 15.120 ;
      LAYER met2 ;
        RECT 56.840 14.560 58.240 14.840 ;
      LAYER met2 ;
        RECT 58.240 14.560 69.440 14.840 ;
      LAYER met2 ;
        RECT 69.440 14.560 70.000 14.840 ;
      LAYER met2 ;
        RECT 70.000 14.560 92.400 14.840 ;
        RECT 56.000 14.000 57.120 14.560 ;
      LAYER met2 ;
        RECT 57.120 14.000 59.080 14.560 ;
      LAYER met2 ;
        RECT 59.080 14.000 92.400 14.560 ;
        RECT 56.000 13.720 56.280 14.000 ;
      LAYER met2 ;
        RECT 56.280 13.720 56.840 14.000 ;
      LAYER met2 ;
        RECT 56.840 13.720 57.120 14.000 ;
      LAYER met2 ;
        RECT 57.120 13.720 57.680 14.000 ;
      LAYER met2 ;
        RECT 57.680 13.720 58.240 14.000 ;
      LAYER met2 ;
        RECT 58.240 13.720 58.800 14.000 ;
      LAYER met2 ;
        RECT 58.800 13.720 92.400 14.000 ;
      LAYER met2 ;
        RECT 55.440 13.440 55.720 13.720 ;
      LAYER met2 ;
        RECT 54.880 13.160 55.160 13.440 ;
      LAYER met2 ;
        RECT 55.160 13.160 55.720 13.440 ;
      LAYER met2 ;
        RECT 50.400 12.880 52.080 13.160 ;
      LAYER met2 ;
        RECT 52.080 12.880 55.720 13.160 ;
      LAYER met2 ;
        RECT 55.720 12.880 56.280 13.720 ;
      LAYER met2 ;
        RECT 56.280 13.440 57.400 13.720 ;
      LAYER met2 ;
        RECT 57.400 13.440 57.960 13.720 ;
      LAYER met2 ;
        RECT 57.960 13.440 58.520 13.720 ;
      LAYER met2 ;
        RECT 58.520 13.440 92.400 13.720 ;
      LAYER met2 ;
        RECT 56.280 12.880 57.120 13.440 ;
      LAYER met2 ;
        RECT 57.120 13.160 57.680 13.440 ;
      LAYER met2 ;
        RECT 57.680 13.160 58.240 13.440 ;
      LAYER met2 ;
        RECT 58.240 13.160 92.400 13.440 ;
        RECT 57.120 12.880 57.400 13.160 ;
      LAYER met2 ;
        RECT 10.920 12.600 11.760 12.880 ;
      LAYER met2 ;
        RECT 11.760 12.600 21.280 12.880 ;
      LAYER met2 ;
        RECT 21.280 12.600 24.360 12.880 ;
      LAYER met2 ;
        RECT 24.360 12.600 26.040 12.880 ;
      LAYER met2 ;
        RECT 26.040 12.600 29.120 12.880 ;
      LAYER met2 ;
        RECT 29.120 12.600 41.720 12.880 ;
      LAYER met2 ;
        RECT 41.720 12.600 45.640 12.880 ;
      LAYER met2 ;
        RECT 45.640 12.600 45.920 12.880 ;
      LAYER met2 ;
        RECT 45.920 12.600 47.600 12.880 ;
      LAYER met2 ;
        RECT 47.600 12.600 49.560 12.880 ;
      LAYER met2 ;
        RECT 49.560 12.600 50.120 12.880 ;
      LAYER met2 ;
        RECT 50.120 12.600 51.240 12.880 ;
      LAYER met2 ;
        RECT 51.240 12.600 55.720 12.880 ;
      LAYER met2 ;
        RECT 55.720 12.600 56.000 12.880 ;
      LAYER met2 ;
        RECT 56.000 12.600 56.840 12.880 ;
      LAYER met2 ;
        RECT 56.840 12.600 57.400 12.880 ;
      LAYER met2 ;
        RECT 57.400 12.600 57.960 13.160 ;
      LAYER met2 ;
        RECT 57.960 12.600 92.400 13.160 ;
      LAYER met2 ;
        RECT 10.920 12.320 11.480 12.600 ;
      LAYER met2 ;
        RECT 11.480 12.320 21.560 12.600 ;
      LAYER met2 ;
        RECT 21.560 12.320 28.840 12.600 ;
      LAYER met2 ;
        RECT 28.840 12.320 42.280 12.600 ;
      LAYER met2 ;
        RECT 42.280 12.320 42.840 12.600 ;
      LAYER met2 ;
        RECT 42.840 12.320 43.400 12.600 ;
      LAYER met2 ;
        RECT 43.400 12.320 43.960 12.600 ;
      LAYER met2 ;
        RECT 43.960 12.320 44.800 12.600 ;
      LAYER met2 ;
        RECT 44.800 12.320 45.360 12.600 ;
      LAYER met2 ;
        RECT 45.360 12.320 46.200 12.600 ;
      LAYER met2 ;
        RECT 46.200 12.320 52.360 12.600 ;
      LAYER met2 ;
        RECT 52.360 12.320 52.640 12.600 ;
      LAYER met2 ;
        RECT 52.640 12.320 56.560 12.600 ;
      LAYER met2 ;
        RECT 56.560 12.320 57.120 12.600 ;
      LAYER met2 ;
        RECT 57.120 12.320 57.680 12.600 ;
      LAYER met2 ;
        RECT 57.680 12.320 92.400 12.600 ;
        RECT 0.000 12.040 4.760 12.320 ;
      LAYER met2 ;
        RECT 4.760 12.040 10.360 12.320 ;
      LAYER met2 ;
        RECT 10.360 12.040 22.120 12.320 ;
      LAYER met2 ;
        RECT 22.120 12.040 28.280 12.320 ;
      LAYER met2 ;
        RECT 28.280 12.040 42.560 12.320 ;
      LAYER met2 ;
        RECT 42.560 12.040 43.120 12.320 ;
      LAYER met2 ;
        RECT 43.120 12.040 46.200 12.320 ;
      LAYER met2 ;
        RECT 46.200 12.040 47.040 12.320 ;
      LAYER met2 ;
        RECT 47.040 12.040 47.600 12.320 ;
        RECT 0.000 11.760 5.320 12.040 ;
      LAYER met2 ;
        RECT 5.320 11.760 10.080 12.040 ;
      LAYER met2 ;
        RECT 10.080 11.760 22.680 12.040 ;
      LAYER met2 ;
        RECT 22.680 11.760 27.720 12.040 ;
      LAYER met2 ;
        RECT 27.720 11.760 42.560 12.040 ;
      LAYER met2 ;
        RECT 42.560 11.760 43.400 12.040 ;
      LAYER met2 ;
        RECT 43.400 11.760 46.480 12.040 ;
      LAYER met2 ;
        RECT 46.480 11.760 47.320 12.040 ;
      LAYER met2 ;
        RECT 47.320 11.760 47.600 12.040 ;
      LAYER met2 ;
        RECT 47.600 11.760 52.080 12.320 ;
      LAYER met2 ;
        RECT 52.080 12.040 52.920 12.320 ;
      LAYER met2 ;
        RECT 52.920 12.040 53.480 12.320 ;
      LAYER met2 ;
        RECT 53.480 12.040 54.040 12.320 ;
      LAYER met2 ;
        RECT 54.040 12.040 54.880 12.320 ;
      LAYER met2 ;
        RECT 54.880 12.040 55.160 12.320 ;
      LAYER met2 ;
        RECT 55.160 12.040 55.720 12.320 ;
      LAYER met2 ;
        RECT 55.720 12.040 56.840 12.320 ;
      LAYER met2 ;
        RECT 56.840 12.040 57.400 12.320 ;
      LAYER met2 ;
        RECT 57.400 12.040 92.400 12.320 ;
        RECT 52.080 11.760 52.640 12.040 ;
      LAYER met2 ;
        RECT 52.640 11.760 53.480 12.040 ;
      LAYER met2 ;
        RECT 53.480 11.760 56.560 12.040 ;
      LAYER met2 ;
        RECT 56.560 11.760 57.120 12.040 ;
      LAYER met2 ;
        RECT 57.120 11.760 92.400 12.040 ;
        RECT 0.000 11.480 6.160 11.760 ;
      LAYER met2 ;
        RECT 6.160 11.480 9.240 11.760 ;
      LAYER met2 ;
        RECT 9.240 11.480 23.800 11.760 ;
      LAYER met2 ;
        RECT 23.800 11.480 26.600 11.760 ;
      LAYER met2 ;
        RECT 26.600 11.480 42.840 11.760 ;
      LAYER met2 ;
        RECT 42.840 11.480 43.680 11.760 ;
      LAYER met2 ;
        RECT 43.680 11.480 46.760 11.760 ;
      LAYER met2 ;
        RECT 46.760 11.480 49.280 11.760 ;
      LAYER met2 ;
        RECT 0.000 11.200 43.120 11.480 ;
      LAYER met2 ;
        RECT 43.120 11.200 43.960 11.480 ;
      LAYER met2 ;
        RECT 43.960 11.200 47.040 11.480 ;
      LAYER met2 ;
        RECT 47.040 11.200 49.280 11.480 ;
      LAYER met2 ;
        RECT 49.280 11.200 49.560 11.760 ;
      LAYER met2 ;
        RECT 49.560 11.480 50.120 11.760 ;
      LAYER met2 ;
        RECT 50.120 11.480 50.680 11.760 ;
      LAYER met2 ;
        RECT 50.680 11.480 52.920 11.760 ;
      LAYER met2 ;
        RECT 52.920 11.480 53.200 11.760 ;
      LAYER met2 ;
        RECT 53.200 11.480 53.480 11.760 ;
      LAYER met2 ;
        RECT 53.480 11.480 56.280 11.760 ;
      LAYER met2 ;
        RECT 56.280 11.480 56.840 11.760 ;
      LAYER met2 ;
        RECT 56.840 11.480 92.400 11.760 ;
      LAYER met2 ;
        RECT 49.560 11.200 50.960 11.480 ;
      LAYER met2 ;
        RECT 0.000 10.920 43.400 11.200 ;
      LAYER met2 ;
        RECT 43.400 10.920 45.080 11.200 ;
      LAYER met2 ;
        RECT 45.080 10.920 47.040 11.200 ;
        RECT 0.000 10.640 43.680 10.920 ;
      LAYER met2 ;
        RECT 43.680 10.640 46.760 10.920 ;
      LAYER met2 ;
        RECT 46.760 10.640 47.040 10.920 ;
      LAYER met2 ;
        RECT 47.040 10.640 50.400 11.200 ;
      LAYER met2 ;
        RECT 50.400 10.640 50.680 11.200 ;
      LAYER met2 ;
        RECT 50.680 10.640 50.960 11.200 ;
      LAYER met2 ;
        RECT 0.000 10.360 45.080 10.640 ;
      LAYER met2 ;
        RECT 45.080 10.360 47.600 10.640 ;
      LAYER met2 ;
        RECT 47.600 10.360 47.880 10.640 ;
        RECT 0.000 9.800 46.480 10.360 ;
      LAYER met2 ;
        RECT 46.480 9.800 47.320 10.360 ;
      LAYER met2 ;
        RECT 47.320 10.080 47.880 10.360 ;
      LAYER met2 ;
        RECT 47.880 10.080 48.440 10.640 ;
      LAYER met2 ;
        RECT 48.440 10.080 49.000 10.640 ;
      LAYER met2 ;
        RECT 49.000 10.360 50.960 10.640 ;
      LAYER met2 ;
        RECT 50.960 10.360 51.240 11.480 ;
      LAYER met2 ;
        RECT 51.240 10.920 52.640 11.480 ;
      LAYER met2 ;
        RECT 52.640 11.200 56.000 11.480 ;
      LAYER met2 ;
        RECT 56.000 11.200 56.560 11.480 ;
      LAYER met2 ;
        RECT 56.560 11.200 92.400 11.480 ;
        RECT 52.640 10.920 54.880 11.200 ;
      LAYER met2 ;
        RECT 54.880 10.920 56.280 11.200 ;
      LAYER met2 ;
        RECT 56.280 10.920 92.400 11.200 ;
      LAYER met2 ;
        RECT 51.240 10.640 52.920 10.920 ;
      LAYER met2 ;
        RECT 52.920 10.640 53.200 10.920 ;
      LAYER met2 ;
        RECT 53.200 10.640 56.000 10.920 ;
      LAYER met2 ;
        RECT 56.000 10.640 92.400 10.920 ;
      LAYER met2 ;
        RECT 51.240 10.360 52.080 10.640 ;
        RECT 49.000 10.080 50.680 10.360 ;
      LAYER met2 ;
        RECT 50.680 10.080 51.520 10.360 ;
      LAYER met2 ;
        RECT 51.520 10.080 52.080 10.360 ;
      LAYER met2 ;
        RECT 52.080 10.080 52.360 10.640 ;
      LAYER met2 ;
        RECT 52.360 10.360 54.880 10.640 ;
      LAYER met2 ;
        RECT 54.880 10.360 92.400 10.640 ;
      LAYER met2 ;
        RECT 52.360 10.080 53.200 10.360 ;
      LAYER met2 ;
        RECT 47.320 9.800 47.600 10.080 ;
      LAYER met2 ;
        RECT 47.600 9.800 48.440 10.080 ;
      LAYER met2 ;
        RECT 48.440 9.800 49.560 10.080 ;
      LAYER met2 ;
        RECT 49.560 9.800 50.120 10.080 ;
      LAYER met2 ;
        RECT 50.120 9.800 51.520 10.080 ;
      LAYER met2 ;
        RECT 51.520 9.800 53.200 10.080 ;
      LAYER met2 ;
        RECT 53.200 9.800 92.400 10.360 ;
        RECT 0.000 9.520 46.760 9.800 ;
        RECT 0.000 9.240 43.400 9.520 ;
      LAYER met2 ;
        RECT 43.400 9.240 44.240 9.520 ;
      LAYER met2 ;
        RECT 44.240 9.240 46.760 9.520 ;
      LAYER met2 ;
        RECT 46.760 9.240 48.160 9.800 ;
      LAYER met2 ;
        RECT 0.000 8.960 42.560 9.240 ;
      LAYER met2 ;
        RECT 42.560 8.960 44.800 9.240 ;
      LAYER met2 ;
        RECT 44.800 8.960 46.480 9.240 ;
      LAYER met2 ;
        RECT 46.480 8.960 48.160 9.240 ;
      LAYER met2 ;
        RECT 48.160 8.960 51.520 9.800 ;
      LAYER met2 ;
        RECT 51.520 9.520 52.920 9.800 ;
      LAYER met2 ;
        RECT 52.920 9.520 92.400 9.800 ;
      LAYER met2 ;
        RECT 51.520 8.960 53.200 9.520 ;
      LAYER met2 ;
        RECT 53.200 9.240 54.880 9.520 ;
      LAYER met2 ;
        RECT 54.880 9.240 56.000 9.520 ;
      LAYER met2 ;
        RECT 56.000 9.240 92.400 9.520 ;
        RECT 53.200 8.960 54.320 9.240 ;
      LAYER met2 ;
        RECT 54.320 8.960 57.120 9.240 ;
      LAYER met2 ;
        RECT 57.120 8.960 92.400 9.240 ;
        RECT 0.000 8.680 41.440 8.960 ;
      LAYER met2 ;
        RECT 41.440 8.680 43.400 8.960 ;
      LAYER met2 ;
        RECT 43.400 8.680 44.240 8.960 ;
      LAYER met2 ;
        RECT 44.240 8.680 45.360 8.960 ;
      LAYER met2 ;
        RECT 45.360 8.680 46.480 8.960 ;
      LAYER met2 ;
        RECT 46.480 8.680 47.880 8.960 ;
      LAYER met2 ;
        RECT 0.000 8.400 40.320 8.680 ;
      LAYER met2 ;
        RECT 40.320 8.400 42.560 8.680 ;
      LAYER met2 ;
        RECT 42.560 8.400 44.800 8.680 ;
      LAYER met2 ;
        RECT 44.800 8.400 45.920 8.680 ;
      LAYER met2 ;
        RECT 45.920 8.400 46.200 8.680 ;
      LAYER met2 ;
        RECT 46.200 8.400 47.040 8.680 ;
      LAYER met2 ;
        RECT 47.040 8.400 47.320 8.680 ;
        RECT 0.000 7.840 39.760 8.400 ;
      LAYER met2 ;
        RECT 39.760 8.120 41.440 8.400 ;
      LAYER met2 ;
        RECT 41.440 8.120 45.360 8.400 ;
      LAYER met2 ;
        RECT 45.360 8.120 46.760 8.400 ;
      LAYER met2 ;
        RECT 46.760 8.120 47.320 8.400 ;
      LAYER met2 ;
        RECT 47.320 8.120 47.880 8.680 ;
      LAYER met2 ;
        RECT 47.880 8.120 51.800 8.960 ;
      LAYER met2 ;
        RECT 51.800 8.680 53.200 8.960 ;
      LAYER met2 ;
        RECT 53.200 8.680 53.760 8.960 ;
      LAYER met2 ;
        RECT 53.760 8.680 54.880 8.960 ;
      LAYER met2 ;
        RECT 54.880 8.680 56.000 8.960 ;
      LAYER met2 ;
        RECT 56.000 8.680 57.960 8.960 ;
      LAYER met2 ;
        RECT 57.960 8.680 92.400 8.960 ;
      LAYER met2 ;
        RECT 39.760 7.840 40.600 8.120 ;
      LAYER met2 ;
        RECT 40.600 7.840 45.920 8.120 ;
        RECT 0.000 7.560 40.040 7.840 ;
      LAYER met2 ;
        RECT 40.040 7.560 41.160 7.840 ;
      LAYER met2 ;
        RECT 41.160 7.560 45.920 7.840 ;
      LAYER met2 ;
        RECT 45.920 7.560 46.760 8.120 ;
      LAYER met2 ;
        RECT 46.760 7.560 47.040 8.120 ;
        RECT 0.000 7.280 40.600 7.560 ;
      LAYER met2 ;
        RECT 40.600 7.280 41.720 7.560 ;
      LAYER met2 ;
        RECT 41.720 7.280 45.920 7.560 ;
      LAYER met2 ;
        RECT 45.920 7.280 46.480 7.560 ;
      LAYER met2 ;
        RECT 46.480 7.280 47.040 7.560 ;
      LAYER met2 ;
        RECT 47.040 7.280 47.600 8.120 ;
      LAYER met2 ;
        RECT 47.600 7.560 51.800 8.120 ;
      LAYER met2 ;
        RECT 51.800 7.840 52.360 8.680 ;
      LAYER met2 ;
        RECT 52.360 8.120 52.640 8.680 ;
      LAYER met2 ;
        RECT 52.640 8.400 54.320 8.680 ;
      LAYER met2 ;
        RECT 54.320 8.400 57.120 8.680 ;
      LAYER met2 ;
        RECT 57.120 8.400 59.080 8.680 ;
      LAYER met2 ;
        RECT 59.080 8.400 92.400 8.680 ;
      LAYER met2 ;
        RECT 52.640 8.120 54.040 8.400 ;
      LAYER met2 ;
        RECT 54.040 8.120 57.960 8.400 ;
      LAYER met2 ;
        RECT 57.960 8.120 59.640 8.400 ;
      LAYER met2 ;
        RECT 52.360 7.840 52.920 8.120 ;
      LAYER met2 ;
        RECT 52.920 7.840 53.480 8.120 ;
      LAYER met2 ;
        RECT 53.480 7.840 58.800 8.120 ;
      LAYER met2 ;
        RECT 58.800 7.840 59.640 8.120 ;
      LAYER met2 ;
        RECT 59.640 7.840 92.400 8.400 ;
      LAYER met2 ;
        RECT 51.800 7.560 52.640 7.840 ;
      LAYER met2 ;
        RECT 47.600 7.280 52.080 7.560 ;
        RECT 0.000 7.000 41.160 7.280 ;
      LAYER met2 ;
        RECT 41.160 7.000 42.280 7.280 ;
      LAYER met2 ;
        RECT 42.280 7.000 45.640 7.280 ;
      LAYER met2 ;
        RECT 45.640 7.000 46.480 7.280 ;
      LAYER met2 ;
        RECT 46.480 7.000 46.760 7.280 ;
        RECT 0.000 6.720 41.720 7.000 ;
      LAYER met2 ;
        RECT 41.720 6.720 42.840 7.000 ;
      LAYER met2 ;
        RECT 42.840 6.720 45.640 7.000 ;
      LAYER met2 ;
        RECT 45.640 6.720 46.200 7.000 ;
      LAYER met2 ;
        RECT 46.200 6.720 46.760 7.000 ;
      LAYER met2 ;
        RECT 46.760 6.720 47.320 7.280 ;
      LAYER met2 ;
        RECT 0.000 6.440 42.280 6.720 ;
      LAYER met2 ;
        RECT 42.280 6.440 43.400 6.720 ;
      LAYER met2 ;
        RECT 43.400 6.440 44.520 6.720 ;
      LAYER met2 ;
        RECT 44.520 6.440 46.200 6.720 ;
      LAYER met2 ;
        RECT 46.200 6.440 46.480 6.720 ;
      LAYER met2 ;
        RECT 46.480 6.440 47.320 6.720 ;
      LAYER met2 ;
        RECT 47.320 6.440 52.080 7.280 ;
      LAYER met2 ;
        RECT 52.080 7.000 52.640 7.560 ;
      LAYER met2 ;
        RECT 52.640 7.280 52.920 7.840 ;
      LAYER met2 ;
        RECT 52.920 7.280 53.760 7.840 ;
      LAYER met2 ;
        RECT 53.760 7.560 58.240 7.840 ;
      LAYER met2 ;
        RECT 58.240 7.560 59.360 7.840 ;
      LAYER met2 ;
        RECT 59.360 7.560 92.400 7.840 ;
        RECT 53.760 7.280 57.680 7.560 ;
      LAYER met2 ;
        RECT 57.680 7.280 58.800 7.560 ;
      LAYER met2 ;
        RECT 58.800 7.280 92.400 7.560 ;
        RECT 52.640 7.000 53.200 7.280 ;
      LAYER met2 ;
        RECT 53.200 7.000 53.760 7.280 ;
      LAYER met2 ;
        RECT 53.760 7.000 57.120 7.280 ;
      LAYER met2 ;
        RECT 57.120 7.000 58.240 7.280 ;
      LAYER met2 ;
        RECT 58.240 7.000 92.400 7.280 ;
        RECT 0.000 6.160 42.840 6.440 ;
      LAYER met2 ;
        RECT 42.840 6.160 47.040 6.440 ;
      LAYER met2 ;
        RECT 0.000 5.880 43.400 6.160 ;
      LAYER met2 ;
        RECT 43.400 5.880 44.520 6.160 ;
      LAYER met2 ;
        RECT 44.520 5.880 45.640 6.160 ;
      LAYER met2 ;
        RECT 45.640 5.880 47.040 6.160 ;
      LAYER met2 ;
        RECT 47.040 5.880 52.080 6.440 ;
      LAYER met2 ;
        RECT 52.080 6.160 52.920 7.000 ;
      LAYER met2 ;
        RECT 52.920 6.160 53.200 7.000 ;
      LAYER met2 ;
        RECT 53.200 6.720 54.040 7.000 ;
      LAYER met2 ;
        RECT 54.040 6.720 56.560 7.000 ;
      LAYER met2 ;
        RECT 56.560 6.720 57.680 7.000 ;
      LAYER met2 ;
        RECT 57.680 6.720 92.400 7.000 ;
      LAYER met2 ;
        RECT 53.200 6.440 54.880 6.720 ;
      LAYER met2 ;
        RECT 54.880 6.440 56.000 6.720 ;
      LAYER met2 ;
        RECT 56.000 6.440 57.120 6.720 ;
      LAYER met2 ;
        RECT 57.120 6.440 92.400 6.720 ;
      LAYER met2 ;
        RECT 53.200 6.160 56.560 6.440 ;
      LAYER met2 ;
        RECT 56.560 6.160 92.400 6.440 ;
      LAYER met2 ;
        RECT 52.080 5.880 54.040 6.160 ;
      LAYER met2 ;
        RECT 54.040 5.880 54.880 6.160 ;
      LAYER met2 ;
        RECT 54.880 5.880 56.000 6.160 ;
      LAYER met2 ;
        RECT 56.000 5.880 92.400 6.160 ;
        RECT 0.000 5.040 46.200 5.880 ;
      LAYER met2 ;
        RECT 46.200 5.600 47.040 5.880 ;
      LAYER met2 ;
        RECT 47.040 5.600 52.360 5.880 ;
      LAYER met2 ;
        RECT 52.360 5.600 54.040 5.880 ;
      LAYER met2 ;
        RECT 54.040 5.600 92.400 5.880 ;
      LAYER met2 ;
        RECT 46.200 5.040 46.760 5.600 ;
      LAYER met2 ;
        RECT 46.760 5.040 52.360 5.600 ;
        RECT 0.000 4.760 45.920 5.040 ;
      LAYER met2 ;
        RECT 45.920 4.760 46.480 5.040 ;
      LAYER met2 ;
        RECT 0.000 4.480 44.800 4.760 ;
      LAYER met2 ;
        RECT 44.800 4.480 46.480 4.760 ;
      LAYER met2 ;
        RECT 0.000 4.200 42.840 4.480 ;
      LAYER met2 ;
        RECT 42.840 4.200 46.480 4.480 ;
      LAYER met2 ;
        RECT 46.480 4.200 52.360 5.040 ;
      LAYER met2 ;
        RECT 52.360 4.760 53.200 5.600 ;
      LAYER met2 ;
        RECT 53.200 4.760 92.400 5.600 ;
      LAYER met2 ;
        RECT 52.360 4.480 54.600 4.760 ;
      LAYER met2 ;
        RECT 54.600 4.480 92.400 4.760 ;
      LAYER met2 ;
        RECT 52.360 4.200 56.560 4.480 ;
      LAYER met2 ;
        RECT 56.560 4.200 92.400 4.480 ;
        RECT 0.000 3.920 42.560 4.200 ;
      LAYER met2 ;
        RECT 42.560 3.920 44.800 4.200 ;
      LAYER met2 ;
        RECT 44.800 3.920 45.640 4.200 ;
      LAYER met2 ;
        RECT 45.640 3.920 46.480 4.200 ;
      LAYER met2 ;
        RECT 46.480 3.920 47.880 4.200 ;
      LAYER met2 ;
        RECT 47.880 3.920 48.160 4.200 ;
      LAYER met2 ;
        RECT 0.000 3.640 42.280 3.920 ;
      LAYER met2 ;
        RECT 42.280 3.640 42.840 3.920 ;
      LAYER met2 ;
        RECT 42.840 3.640 45.640 3.920 ;
      LAYER met2 ;
        RECT 45.640 3.640 46.760 3.920 ;
      LAYER met2 ;
        RECT 46.760 3.640 47.600 3.920 ;
      LAYER met2 ;
        RECT 47.600 3.640 48.160 3.920 ;
      LAYER met2 ;
        RECT 48.160 3.640 49.280 4.200 ;
      LAYER met2 ;
        RECT 49.280 3.920 49.560 4.200 ;
      LAYER met2 ;
        RECT 49.560 3.920 50.960 4.200 ;
      LAYER met2 ;
        RECT 50.960 3.920 51.240 4.200 ;
      LAYER met2 ;
        RECT 51.240 3.920 52.360 4.200 ;
      LAYER met2 ;
        RECT 52.360 3.920 53.200 4.200 ;
      LAYER met2 ;
        RECT 53.200 3.920 54.600 4.200 ;
      LAYER met2 ;
        RECT 54.600 3.920 56.840 4.200 ;
      LAYER met2 ;
        RECT 56.840 3.920 92.400 4.200 ;
      LAYER met2 ;
        RECT 49.280 3.640 49.840 3.920 ;
      LAYER met2 ;
        RECT 0.000 3.360 42.000 3.640 ;
      LAYER met2 ;
        RECT 42.000 3.360 42.560 3.640 ;
      LAYER met2 ;
        RECT 0.000 3.080 41.720 3.360 ;
      LAYER met2 ;
        RECT 41.720 3.080 42.560 3.360 ;
      LAYER met2 ;
        RECT 42.560 3.080 45.360 3.640 ;
        RECT 0.000 2.520 41.440 3.080 ;
      LAYER met2 ;
        RECT 41.440 2.800 42.280 3.080 ;
      LAYER met2 ;
        RECT 42.280 2.800 45.360 3.080 ;
      LAYER met2 ;
        RECT 45.360 2.800 45.920 3.640 ;
      LAYER met2 ;
        RECT 45.920 3.360 46.200 3.640 ;
      LAYER met2 ;
        RECT 46.200 3.360 46.760 3.640 ;
      LAYER met2 ;
        RECT 46.760 3.360 47.320 3.640 ;
      LAYER met2 ;
        RECT 47.320 3.360 48.160 3.640 ;
      LAYER met2 ;
        RECT 48.160 3.360 49.000 3.640 ;
      LAYER met2 ;
        RECT 49.000 3.360 49.840 3.640 ;
      LAYER met2 ;
        RECT 49.840 3.360 50.960 3.920 ;
      LAYER met2 ;
        RECT 50.960 3.640 51.520 3.920 ;
      LAYER met2 ;
        RECT 51.520 3.640 52.640 3.920 ;
      LAYER met2 ;
        RECT 52.640 3.640 53.200 3.920 ;
      LAYER met2 ;
        RECT 53.200 3.640 56.280 3.920 ;
      LAYER met2 ;
        RECT 56.280 3.640 57.120 3.920 ;
      LAYER met2 ;
        RECT 57.120 3.640 92.400 3.920 ;
      LAYER met2 ;
        RECT 50.960 3.360 51.800 3.640 ;
      LAYER met2 ;
        RECT 51.800 3.360 52.640 3.640 ;
      LAYER met2 ;
        RECT 52.640 3.360 53.480 3.640 ;
      LAYER met2 ;
        RECT 53.480 3.360 56.560 3.640 ;
      LAYER met2 ;
        RECT 56.560 3.360 57.400 3.640 ;
      LAYER met2 ;
        RECT 57.400 3.360 92.400 3.640 ;
        RECT 45.920 2.800 46.480 3.360 ;
      LAYER met2 ;
        RECT 46.480 2.800 47.600 3.360 ;
      LAYER met2 ;
        RECT 47.600 3.080 47.880 3.360 ;
      LAYER met2 ;
        RECT 47.880 3.080 48.440 3.360 ;
      LAYER met2 ;
        RECT 48.440 3.080 49.000 3.360 ;
      LAYER met2 ;
        RECT 49.000 3.080 49.280 3.360 ;
      LAYER met2 ;
        RECT 49.280 3.080 49.560 3.360 ;
      LAYER met2 ;
        RECT 49.560 3.080 50.120 3.360 ;
      LAYER met2 ;
        RECT 47.600 2.800 48.160 3.080 ;
      LAYER met2 ;
        RECT 48.160 2.800 48.440 3.080 ;
      LAYER met2 ;
        RECT 48.440 2.800 48.720 3.080 ;
      LAYER met2 ;
        RECT 48.720 2.800 49.280 3.080 ;
      LAYER met2 ;
        RECT 49.280 2.800 49.840 3.080 ;
      LAYER met2 ;
        RECT 49.840 2.800 50.120 3.080 ;
      LAYER met2 ;
        RECT 50.120 2.800 50.680 3.360 ;
      LAYER met2 ;
        RECT 50.680 3.080 51.240 3.360 ;
      LAYER met2 ;
        RECT 51.240 3.080 51.520 3.360 ;
      LAYER met2 ;
        RECT 51.520 3.080 51.800 3.360 ;
      LAYER met2 ;
        RECT 51.800 3.080 52.360 3.360 ;
      LAYER met2 ;
        RECT 52.360 3.080 53.480 3.360 ;
      LAYER met2 ;
        RECT 53.480 3.080 56.840 3.360 ;
      LAYER met2 ;
        RECT 56.840 3.080 57.680 3.360 ;
        RECT 50.680 2.800 50.960 3.080 ;
      LAYER met2 ;
        RECT 50.960 2.800 51.520 3.080 ;
      LAYER met2 ;
        RECT 51.520 2.800 52.080 3.080 ;
      LAYER met2 ;
        RECT 52.080 2.800 52.360 3.080 ;
      LAYER met2 ;
        RECT 52.360 2.800 53.760 3.080 ;
      LAYER met2 ;
        RECT 53.760 2.800 57.120 3.080 ;
      LAYER met2 ;
        RECT 57.120 2.800 57.680 3.080 ;
      LAYER met2 ;
        RECT 57.680 2.800 92.400 3.360 ;
      LAYER met2 ;
        RECT 41.440 2.520 42.000 2.800 ;
      LAYER met2 ;
        RECT 42.000 2.520 45.360 2.800 ;
      LAYER met2 ;
        RECT 45.360 2.520 46.200 2.800 ;
      LAYER met2 ;
        RECT 46.200 2.520 46.760 2.800 ;
      LAYER met2 ;
        RECT 46.760 2.520 47.320 2.800 ;
      LAYER met2 ;
        RECT 0.000 2.240 41.160 2.520 ;
      LAYER met2 ;
        RECT 41.160 2.240 41.720 2.520 ;
      LAYER met2 ;
        RECT 41.720 2.240 45.080 2.520 ;
      LAYER met2 ;
        RECT 45.080 2.240 47.320 2.520 ;
      LAYER met2 ;
        RECT 47.320 2.240 48.160 2.800 ;
      LAYER met2 ;
        RECT 48.160 2.240 49.000 2.800 ;
      LAYER met2 ;
        RECT 49.000 2.520 49.840 2.800 ;
      LAYER met2 ;
        RECT 49.840 2.520 50.960 2.800 ;
      LAYER met2 ;
        RECT 50.960 2.520 51.800 2.800 ;
      LAYER met2 ;
        RECT 51.800 2.520 54.040 2.800 ;
      LAYER met2 ;
        RECT 54.040 2.520 57.400 2.800 ;
      LAYER met2 ;
        RECT 57.400 2.520 57.960 2.800 ;
      LAYER met2 ;
        RECT 57.960 2.520 92.400 2.800 ;
        RECT 49.000 2.240 50.120 2.520 ;
      LAYER met2 ;
        RECT 50.120 2.240 50.680 2.520 ;
      LAYER met2 ;
        RECT 50.680 2.240 51.800 2.520 ;
      LAYER met2 ;
        RECT 51.800 2.240 53.480 2.520 ;
      LAYER met2 ;
        RECT 53.480 2.240 53.760 2.520 ;
      LAYER met2 ;
        RECT 53.760 2.240 54.320 2.520 ;
      LAYER met2 ;
        RECT 54.320 2.240 57.680 2.520 ;
      LAYER met2 ;
        RECT 57.680 2.240 58.240 2.520 ;
      LAYER met2 ;
        RECT 58.240 2.240 92.400 2.520 ;
        RECT 0.000 1.960 40.880 2.240 ;
      LAYER met2 ;
        RECT 40.880 1.960 41.440 2.240 ;
      LAYER met2 ;
        RECT 41.440 1.960 44.800 2.240 ;
      LAYER met2 ;
        RECT 44.800 1.960 45.360 2.240 ;
      LAYER met2 ;
        RECT 45.360 1.960 45.920 2.240 ;
      LAYER met2 ;
        RECT 45.920 1.960 53.480 2.240 ;
      LAYER met2 ;
        RECT 53.480 1.960 54.040 2.240 ;
      LAYER met2 ;
        RECT 54.040 1.960 54.600 2.240 ;
      LAYER met2 ;
        RECT 54.600 1.960 57.960 2.240 ;
      LAYER met2 ;
        RECT 57.960 1.960 58.520 2.240 ;
      LAYER met2 ;
        RECT 58.520 1.960 92.400 2.240 ;
        RECT 0.000 1.680 40.600 1.960 ;
      LAYER met2 ;
        RECT 40.600 1.680 41.160 1.960 ;
      LAYER met2 ;
        RECT 41.160 1.680 44.520 1.960 ;
      LAYER met2 ;
        RECT 44.520 1.680 45.080 1.960 ;
      LAYER met2 ;
        RECT 45.080 1.680 45.920 1.960 ;
      LAYER met2 ;
        RECT 45.920 1.680 53.200 1.960 ;
      LAYER met2 ;
        RECT 53.200 1.680 54.320 1.960 ;
      LAYER met2 ;
        RECT 54.320 1.680 54.880 1.960 ;
      LAYER met2 ;
        RECT 54.880 1.680 58.240 1.960 ;
      LAYER met2 ;
        RECT 58.240 1.680 58.800 1.960 ;
      LAYER met2 ;
        RECT 58.800 1.680 92.400 1.960 ;
        RECT 0.000 1.400 40.320 1.680 ;
      LAYER met2 ;
        RECT 40.320 1.400 40.880 1.680 ;
      LAYER met2 ;
        RECT 40.880 1.400 43.400 1.680 ;
      LAYER met2 ;
        RECT 43.400 1.400 44.800 1.680 ;
      LAYER met2 ;
        RECT 44.800 1.400 45.920 1.680 ;
      LAYER met2 ;
        RECT 45.920 1.400 46.760 1.680 ;
      LAYER met2 ;
        RECT 46.760 1.400 47.320 1.680 ;
      LAYER met2 ;
        RECT 47.320 1.400 47.880 1.680 ;
      LAYER met2 ;
        RECT 0.000 1.120 40.040 1.400 ;
      LAYER met2 ;
        RECT 40.040 1.120 40.600 1.400 ;
      LAYER met2 ;
        RECT 40.600 1.120 41.160 1.400 ;
      LAYER met2 ;
        RECT 41.160 1.120 44.520 1.400 ;
      LAYER met2 ;
        RECT 44.520 1.120 45.920 1.400 ;
      LAYER met2 ;
        RECT 45.920 1.120 47.880 1.400 ;
      LAYER met2 ;
        RECT 47.880 1.120 50.680 1.680 ;
      LAYER met2 ;
        RECT 50.680 1.400 51.520 1.680 ;
      LAYER met2 ;
        RECT 51.520 1.400 52.080 1.680 ;
      LAYER met2 ;
        RECT 52.080 1.400 52.920 1.680 ;
      LAYER met2 ;
        RECT 52.920 1.400 54.600 1.680 ;
      LAYER met2 ;
        RECT 54.600 1.400 56.000 1.680 ;
      LAYER met2 ;
        RECT 56.000 1.400 58.520 1.680 ;
      LAYER met2 ;
        RECT 58.520 1.400 59.080 1.680 ;
      LAYER met2 ;
        RECT 59.080 1.400 92.400 1.680 ;
      LAYER met2 ;
        RECT 50.680 1.120 52.640 1.400 ;
      LAYER met2 ;
        RECT 52.640 1.120 54.880 1.400 ;
      LAYER met2 ;
        RECT 54.880 1.120 57.960 1.400 ;
      LAYER met2 ;
        RECT 57.960 1.120 58.800 1.400 ;
      LAYER met2 ;
        RECT 58.800 1.120 59.360 1.400 ;
      LAYER met2 ;
        RECT 59.360 1.120 92.400 1.400 ;
        RECT 0.000 0.560 39.760 1.120 ;
      LAYER met2 ;
        RECT 39.760 0.840 43.400 1.120 ;
      LAYER met2 ;
        RECT 43.400 0.840 46.200 1.120 ;
      LAYER met2 ;
        RECT 46.200 0.840 47.600 1.120 ;
      LAYER met2 ;
        RECT 47.600 0.840 50.960 1.120 ;
      LAYER met2 ;
        RECT 50.960 0.840 52.640 1.120 ;
      LAYER met2 ;
        RECT 52.640 0.840 56.000 1.120 ;
      LAYER met2 ;
        RECT 56.000 0.840 59.640 1.120 ;
        RECT 39.760 0.560 41.160 0.840 ;
      LAYER met2 ;
        RECT 41.160 0.560 51.240 0.840 ;
      LAYER met2 ;
        RECT 51.240 0.560 52.080 0.840 ;
      LAYER met2 ;
        RECT 52.080 0.560 57.960 0.840 ;
      LAYER met2 ;
        RECT 57.960 0.560 59.640 0.840 ;
      LAYER met2 ;
        RECT 59.640 0.560 92.400 1.120 ;
        RECT 0.000 0.000 92.400 0.560 ;
      LAYER met3 ;
        RECT 0.000 0.000 92.400 29.400 ;
      LAYER met4 ;
        RECT 0.000 0.000 92.400 29.400 ;
      LAYER met5 ;
        RECT 0.000 0.000 92.400 29.400 ;
  END
END tt09ball4_logo
END LIBRARY

