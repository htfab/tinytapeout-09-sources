magic
tech sky130A
magscale 1 2
timestamp 1730926491
<< locali >>
rect -2020 940 -1060 1040
rect -1660 880 -1400 940
rect -1840 460 -1740 640
rect -1520 460 -1420 640
rect -1940 -320 -1840 -140
rect -1640 -320 -1540 -140
rect -1520 -320 -1420 -140
rect -1220 -320 -1120 -140
rect -1660 -620 -1400 -560
rect -2020 -720 -1060 -620
<< metal1 >>
rect -2020 740 -1640 840
rect -1580 740 -1320 840
rect -2020 220 -1920 740
rect -1580 600 -1480 740
rect -1640 500 -1480 600
rect -1320 500 -1060 600
rect -1580 380 -1480 500
rect -1740 220 -1640 380
rect -2020 120 -1640 220
rect -2020 -420 -1920 120
rect -1740 -40 -1640 120
rect -1580 280 -1320 380
rect -1580 60 -1480 280
rect -1580 -40 -1220 60
rect -1780 -200 -1700 -180
rect -1780 -260 -1760 -200
rect -1780 -280 -1700 -260
rect -1580 -200 -1480 -40
rect -1580 -260 -1560 -200
rect -1500 -260 -1480 -200
rect -1580 -420 -1480 -260
rect -1360 -200 -1280 -180
rect -1360 -260 -1340 -200
rect -1360 -280 -1280 -260
rect -1160 -200 -1060 500
rect -1160 -260 -1140 -200
rect -1080 -260 -1060 -200
rect -1160 -280 -1060 -260
rect -2020 -520 -1740 -420
rect -1580 -520 -1320 -420
<< via1 >>
rect -1760 -260 -1700 -200
rect -1560 -260 -1500 -200
rect -1340 -260 -1280 -200
rect -1140 -260 -1080 -200
<< metal2 >>
rect -1780 -200 -1480 -180
rect -1780 -260 -1760 -200
rect -1700 -260 -1560 -200
rect -1500 -260 -1480 -200
rect -1780 -280 -1480 -260
rect -1360 -200 -1060 -180
rect -1360 -260 -1340 -200
rect -1280 -260 -1140 -200
rect -1080 -260 -1060 -200
rect -1360 -280 -1060 -260
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_0
timestamp 1730922800
transform 1 0 -1689 0 1 560
box -211 -360 211 360
use sky130_fd_pr__nfet_01v8_NRQ53D  sky130_fd_pr__nfet_01v8_NRQ53D_2
timestamp 1730922800
transform 1 0 -1373 0 1 560
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_0
timestamp 1730925979
transform 1 0 -1317 0 1 -231
box -263 -369 263 369
use sky130_fd_pr__pfet_01v8_XJBLHL  sky130_fd_pr__pfet_01v8_XJBLHL_2
timestamp 1730925979
transform 1 0 -1737 0 1 -231
box -263 -369 263 369
<< labels >>
rlabel locali -2020 -720 -1920 -620 1 VPWR
port 1 n
rlabel locali -2020 940 -1920 1040 1 VGND
port 2 n
rlabel metal1 -2020 120 -1920 220 1 IN
port 3 n
rlabel metal1 -1160 120 -1060 220 1 Q_P
port 4 n
rlabel metal1 -1580 120 -1480 220 1 Q_N
port 5 n
<< end >>
