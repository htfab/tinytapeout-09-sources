*SWTCH_GATE_SKY130NM/SWTCH_GATE
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SWTCH_GATE_lpe.spi
#else
.include ../../../work/xsch/SWTCH_GATE.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VGND VGND GND dc 0
VPWR VPWR GND pwl 0 0 100p {AVDD}

VP CTRL_P GND pwl 0 0 100p {AVDD}
VN CTRL_N GND pwl 0 0 100p 0

VX X GND pwl 0 0 100p {AVDD}

IY Y GND pwl 0 0 1n 0 2n 100u

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VPWR VGND CTRL_P CTRL_N X Y SWTCH_GATE

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.probe v(VPWR) v(VGND) v(CTRL_P) v(CTRL_N) v(X) v(Y)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 10n 1p
write
quit
#endif

.endc

.end
