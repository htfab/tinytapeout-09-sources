* NGSPICE file created from saff_2_parax.ext - technology: sky130A

.subckt saff_2_parax clk q nq VSS1 VDD2 VSS2 nd d VDD1
X0 VSS2.t26 clk.t0 a_570_510.t8 VSS2.t25 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X1 nq.t3 sense_amplifier_0.out2.t4 a_1336_n1386# VSS2.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X2 a_570_510.t2 d.t0 a_658_510# VSS2.t2 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X3 VSS2.t24 clk.t1 a_570_510.t9 VSS2.t23 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4 q.t1 a_690_n1522# VSS2.t9 VSS2.t8 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X5 a_958_n1386# sense_amplifier_0.out1.t4 q.t2 VSS2.t11 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X6 a_834_510.t3 sense_amplifier_0.out1.t5 sense_amplifier_0.out2.t1 VSS2.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X7 VDD1.t5 clk.t2 sense_amplifier_0.out2.t2 VDD1.t4 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X8 a_658_510# d.t1 a_570_510.t1 VSS2.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X9 sense_amplifier_0.out1.t0 clk.t3 VDD1.t3 VDD1.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X10 a_570_510.t12 nd.t0 a_834_510.t5 VSS2.t10 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X11 VDD2.t13 sense_amplifier_0.out2.t5 nq.t2 VDD2.t12 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X12 sense_amplifier_0.out1.t3 sense_amplifier_0.out2.t6 a_658_510# VSS2.t13 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X13 VDD2.t1 nq.t4 a_958_n952# VDD2.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X14 a_658_510# d.t2 a_570_510.t5 VSS2.t16 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X15 VSS2.t29 sense_amplifier_0.out2.t7 a_690_n1522# VSS2.t28 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X16 a_834_510.t0 nd.t1 a_570_510.t0 VSS2.t1 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X17 a_570_510.t10 clk.t4 VSS2.t22 VSS2.t21 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X18 a_570_510.t11 clk.t5 VSS2.t20 VSS2.t19 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X19 q.t3 sense_amplifier_0.out1.t6 VDD2.t6 VDD2.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X20 a_1374_n306# sense_amplifier_0.out1.t7 VSS2.t31 VSS2.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X21 sense_amplifier_0.out2.t3 sense_amplifier_0.out1.t8 VDD1.t1 VDD1.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X22 a_1336_n1386# q.t4 VSS2.t4 VSS2.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X23 a_834_510.t4 nd.t2 a_570_510.t6 VSS2.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X24 VSS2.t15 nq.t5 a_958_n1386# VSS2.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X25 sense_amplifier_0.out2.t0 sense_amplifier_0.out1.t9 a_834_510.t2 VSS2.t10 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X26 a_570_510.t3 nd.t3 a_834_510.t1 VSS2.t5 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X27 nq.t1 a_1374_n306# a_1336_n952# VDD2.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X28 a_658_510# sense_amplifier_0.out2.t8 sense_amplifier_0.out1.t2 VSS2.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X29 a_570_510.t4 d.t3 a_658_510# VSS2.t13 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X30 a_958_n952# a_690_n1522# q.t0 VDD2.t9 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X31 VSS2.t7 a_1374_n306# nq.t0 VSS2.t6 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X32 VDD1.t7 sense_amplifier_0.out2.t9 sense_amplifier_0.out1.t1 VDD1.t6 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X33 VSS2.t18 clk.t6 a_570_510.t7 VSS2.t17 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X34 a_1374_n306# sense_amplifier_0.out1.t10 VDD2.t4 VDD2.t3 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X35 a_1336_n952# q.t5 VDD2.t8 VDD2.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X36 VDD2.t11 sense_amplifier_0.out2.t10 a_690_n1522# VDD2.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
R0 clk.n0 clk.t3 851.506
R1 clk.n0 clk.t2 850.414
R2 clk.n1 clk.t6 665.16
R3 clk.n1 clk.t5 523.774
R4 clk.n2 clk.t1 523.774
R5 clk.n3 clk.t4 523.774
R6 clk.n4 clk.t0 523.774
R7 clk.n5 clk.n4 213.51
R8 clk.n4 clk.n3 141.387
R9 clk.n3 clk.n2 141.387
R10 clk.n2 clk.n1 141.387
R11 clk clk.n5 11.8482
R12 clk.n5 clk.n0 1.05649
R13 a_570_510.n9 a_570_510.t1 32.0282
R14 a_570_510.n4 a_570_510.n3 25.7663
R15 a_570_510.n7 a_570_510.n1 25.75
R16 a_570_510.n8 a_570_510.n0 25.75
R17 a_570_510.n10 a_570_510.n9 25.75
R18 a_570_510.n4 a_570_510.n2 25.288
R19 a_570_510.n6 a_570_510.n5 24.288
R20 a_570_510.n5 a_570_510.t7 5.8005
R21 a_570_510.n5 a_570_510.t12 5.8005
R22 a_570_510.n2 a_570_510.t9 5.8005
R23 a_570_510.n2 a_570_510.t11 5.8005
R24 a_570_510.n3 a_570_510.t8 5.8005
R25 a_570_510.n3 a_570_510.t10 5.8005
R26 a_570_510.n1 a_570_510.t6 5.8005
R27 a_570_510.n1 a_570_510.t2 5.8005
R28 a_570_510.n0 a_570_510.t5 5.8005
R29 a_570_510.n0 a_570_510.t3 5.8005
R30 a_570_510.t0 a_570_510.n10 5.8005
R31 a_570_510.n10 a_570_510.t4 5.8005
R32 a_570_510.n7 a_570_510.n6 1.94072
R33 a_570_510.n6 a_570_510.n4 1.47876
R34 a_570_510.n8 a_570_510.n7 0.478761
R35 a_570_510.n9 a_570_510.n8 0.478761
R36 VSS2.n47 VSS2.n46 37135.8
R37 VSS2.n46 VSS2.n10 11686.1
R38 VSS2.n49 VSS2.n47 10321.3
R39 VSS2.n39 VSS2.n22 4042.48
R40 VSS2.n32 VSS2.n22 3140.17
R41 VSS2.n40 VSS2.n12 3120.05
R42 VSS2.n44 VSS2.n12 2350.81
R43 VSS2.n53 VSS2.n7 2235.89
R44 VSS2.n48 VSS2.n8 2230.09
R45 VSS2.n37 VSS2.n22 1915.82
R46 VSS2.n38 VSS2.n37 1832.1
R47 VSS2.n44 VSS2.n11 1562.99
R48 VSS2.n50 VSS2.n8 1411.83
R49 VSS2.n26 VSS2.n23 1226.74
R50 VSS2.n39 VSS2.n38 1068.72
R51 VSS2.n10 VSS2.t30 994.611
R52 VSS2.n51 VSS2.t14 955.091
R53 VSS2.t28 VSS2.n49 955.091
R54 VSS2.n52 VSS2.t3 935.33
R55 VSS2.n32 VSS2.n26 742.855
R56 VSS2.t30 VSS2.t6 579.641
R57 VSS2.t6 VSS2.t27 579.641
R58 VSS2.t27 VSS2.t3 579.641
R59 VSS2.t14 VSS2.t11 579.641
R60 VSS2.t11 VSS2.t8 579.641
R61 VSS2.t8 VSS2.t28 579.641
R62 VSS2.n47 VSS2.n9 392.099
R63 VSS2.n26 VSS2.n11 356.277
R64 VSS2.n45 VSS2.t25 338.017
R65 VSS2.t0 VSS2.n9 338.017
R66 VSS2.n40 VSS2.n39 281.135
R67 VSS2.n27 VSS2.n20 262.659
R68 VSS2.n31 VSS2.n27 204.031
R69 VSS2.n42 VSS2.n41 202.725
R70 VSS2.t23 VSS2.t21 169.975
R71 VSS2.t17 VSS2.t19 169.975
R72 VSS2.t10 VSS2.t17 169.975
R73 VSS2.t12 VSS2.t10 169.975
R74 VSS2.t2 VSS2.t12 169.975
R75 VSS2.t16 VSS2.t2 169.975
R76 VSS2.t5 VSS2.t1 169.975
R77 VSS2.t1 VSS2.t13 169.975
R78 VSS2.t13 VSS2.t0 169.975
R79 VSS2.n33 VSS2.t23 168.042
R80 VSS2.n43 VSS2.n42 152.744
R81 VSS2.n55 VSS2.n6 138.52
R82 VSS2.n54 VSS2.n0 138.144
R83 VSS2.n27 VSS2.n24 124.481
R84 VSS2.n28 VSS2.n24 119.04
R85 VSS2.n13 VSS2.n11 117.001
R86 VSS2.n25 VSS2.n11 117.001
R87 VSS2.n7 VSS2.n6 104.257
R88 VSS2.n48 VSS2.n0 104.257
R89 VSS2.n43 VSS2.n13 101.555
R90 VSS2.n10 VSS2.n7 97.5005
R91 VSS2.n49 VSS2.n48 97.5005
R92 VSS2.n50 VSS2.n2 92.3255
R93 VSS2.n25 VSS2.t25 86.9189
R94 VSS2.n3 VSS2.t4 84.5161
R95 VSS2.n58 VSS2.t15 84.5161
R96 VSS2.t21 VSS2.n25 83.0558
R97 VSS2.n36 VSS2.t5 83.0558
R98 VSS2.n30 VSS2.n29 79.7072
R99 VSS2.n32 VSS2.n31 73.1255
R100 VSS2.n33 VSS2.n32 73.1255
R101 VSS2.n51 VSS2.n50 73.1255
R102 VSS2.n54 VSS2.n2 72.5338
R103 VSS2.n28 VSS2.n20 69.4405
R104 VSS2.n5 VSS2.n4 67.1161
R105 VSS2.n59 VSS2.n1 67.1161
R106 VSS2.n34 VSS2.t16 59.8776
R107 VSS2.n37 VSS2.n24 53.1823
R108 VSS2.n37 VSS2.n36 53.1823
R109 VSS2.n29 VSS2.n23 48.7505
R110 VSS2.n34 VSS2.n23 48.7505
R111 VSS2.n31 VSS2.n30 48.2672
R112 VSS2.n27 VSS2.n22 45.0005
R113 VSS2.n35 VSS2.n22 45.0005
R114 VSS2.n44 VSS2.n43 39.0005
R115 VSS2.n45 VSS2.n44 39.0005
R116 VSS2.n38 VSS2.n23 34.4755
R117 VSS2.n14 VSS2.t26 31.7728
R118 VSS2.n17 VSS2.n16 25.9728
R119 VSS2.n18 VSS2.n15 25.9728
R120 VSS2.n35 VSS2.n34 23.1787
R121 VSS2.n30 VSS2.n13 23.1494
R122 VSS2.n41 VSS2.n40 22.5005
R123 VSS2.n40 VSS2.n9 22.5005
R124 VSS2.n52 VSS2.n51 19.761
R125 VSS2.n46 VSS2.n45 19.3157
R126 VSS2.n41 VSS2.n20 18.2672
R127 VSS2.n4 VSS2.t31 17.4005
R128 VSS2.n4 VSS2.t7 17.4005
R129 VSS2.n1 VSS2.t9 17.4005
R130 VSS2.n1 VSS2.t29 17.4005
R131 VSS2.n55 VSS2.n53 17.2064
R132 VSS2.n53 VSS2.n52 17.2064
R133 VSS2.n42 VSS2.n12 15.3952
R134 VSS2.t12 VSS2.n12 15.3952
R135 VSS2.n16 VSS2.t22 5.8005
R136 VSS2.n16 VSS2.t24 5.8005
R137 VSS2.n15 VSS2.t20 5.8005
R138 VSS2.n15 VSS2.t18 5.8005
R139 VSS2.n53 VSS2.n8 5.79462
R140 VSS2.n36 VSS2.n35 3.86354
R141 VSS2.n6 VSS2.n5 2.60207
R142 VSS2.n57 VSS2.n2 2.39175
R143 VSS2.n60 VSS2.n0 2.3631
R144 VSS2.n29 VSS2.n28 2.2405
R145 VSS2.t19 VSS2.n33 1.93202
R146 VSS2.n41 VSS2.n21 1.56378
R147 VSS2.n43 VSS2.n14 1.51802
R148 VSS2.n21 VSS2.n19 0.785098
R149 VSS2.n56 VSS2.n55 0.58175
R150 VSS2.n21 VSS1 0.522821
R151 VSS2.n42 VSS2.n19 0.517167
R152 VSS2.n55 VSS2.n54 0.376971
R153 VSS2.n5 VSS2.n3 0.324029
R154 VSS2.n59 VSS2.n58 0.324029
R155 VSS2.n19 VSS2.n18 0.246036
R156 VSS2.n60 VSS2.n59 0.232118
R157 VSS2.n17 VSS2.n14 0.196929
R158 VSS2.n18 VSS2.n17 0.196929
R159 VSS2.n58 VSS2.n57 0.124275
R160 VSS2.n56 VSS2.n3 0.120598
R161 VSS2 VSS2.n60 0.113245
R162 VSS2.n57 VSS2.n56 0.00417647
R163 sense_amplifier_0.out2.n1 sense_amplifier_0.out2.t9 879.481
R164 sense_amplifier_0.out2.n4 sense_amplifier_0.out2.t10 742.783
R165 sense_amplifier_0.out2.n5 sense_amplifier_0.out2.t8 665.16
R166 sense_amplifier_0.out2.n2 sense_amplifier_0.out2.t5 623.388
R167 sense_amplifier_0.out2.n5 sense_amplifier_0.out2.t6 523.774
R168 sense_amplifier_0.out2.n2 sense_amplifier_0.out2.t4 431.807
R169 sense_amplifier_0.out2.n4 sense_amplifier_0.out2.t7 427.875
R170 sense_amplifier_0.out2.n1 sense_amplifier_0.out2.n5 357.26
R171 sense_amplifier_0.out2 sense_amplifier_0.out2.n2 208.537
R172 sense_amplifier_0.out2 sense_amplifier_0.out2.n4 168.077
R173 sense_amplifier_0.out2.n0 sense_amplifier_0.out2.n3 75.5326
R174 sense_amplifier_0.out2.n0 sense_amplifier_0.out2.t1 31.2347
R175 sense_amplifier_0.out2.n6 sense_amplifier_0.out2.t0 31.2347
R176 sense_amplifier_0.out2.n1 sense_amplifier_0.out2 11.1806
R177 sense_amplifier_0.out2 sense_amplifier_0.out2.n6 10.5958
R178 sense_amplifier_0.out2.n3 sense_amplifier_0.out2.t2 9.52217
R179 sense_amplifier_0.out2.n3 sense_amplifier_0.out2.t3 9.52217
R180 sense_amplifier_0.out2.n0 sense_amplifier_0.out2.n1 0.803118
R181 sense_amplifier_0.out2.n6 sense_amplifier_0.out2.n0 0.478761
R182 nq.n1 nq.t4 567.446
R183 nq.n1 nq.t5 400.353
R184 nq.n2 nq.n1 162.399
R185 nq.n2 nq.n0 75.2282
R186 nq.n4 nq.n3 66.3172
R187 nq.n3 nq.t0 17.4005
R188 nq.n3 nq.t3 17.4005
R189 nq.n0 nq.t2 9.52217
R190 nq.n0 nq.t1 9.52217
R191 nq nq.n4 5.09289
R192 nq.n4 nq.n2 0.658109
R193 d.n1 d.t3 572.12
R194 d.n1 d.t1 572.12
R195 d.n0 d.t0 572.12
R196 d.n0 d.t2 572.12
R197 d.n2 d.n0 166.468
R198 d.n2 d.n1 165.8
R199 d d.n2 16.0275
R200 q.n1 q.t5 734.539
R201 q.n1 q.t4 233.26
R202 q.n2 q.n1 162.399
R203 q.n2 q.n0 75.5108
R204 q.n4 q.n3 66.3172
R205 q.n3 q.t2 17.4005
R206 q.n3 q.t1 17.4005
R207 q.n0 q.t0 9.52217
R208 q.n0 q.t3 9.52217
R209 q q.n4 5.08746
R210 q.n4 q.n2 0.3755
R211 sense_amplifier_0.out1.n6 sense_amplifier_0.out1.t8 890.727
R212 sense_amplifier_0.out1.n0 sense_amplifier_0.out1.t10 742.783
R213 sense_amplifier_0.out1.n7 sense_amplifier_0.out1.t9 665.16
R214 sense_amplifier_0.out1.n2 sense_amplifier_0.out1.t6 623.388
R215 sense_amplifier_0.out1.n7 sense_amplifier_0.out1.t5 523.774
R216 sense_amplifier_0.out1.n2 sense_amplifier_0.out1.t4 431.807
R217 sense_amplifier_0.out1.n0 sense_amplifier_0.out1.t7 427.875
R218 sense_amplifier_0.out1.n8 sense_amplifier_0.out1.n7 364.733
R219 sense_amplifier_0.out1 sense_amplifier_0.out1.n2 208.5
R220 sense_amplifier_0.out1 sense_amplifier_0.out1.n0 168.007
R221 sense_amplifier_0.out1.n5 sense_amplifier_0.out1.n1 75.2663
R222 sense_amplifier_0.out1.n4 sense_amplifier_0.out1.t3 31.2728
R223 sense_amplifier_0.out1.n3 sense_amplifier_0.out1.t2 31.0337
R224 sense_amplifier_0.out1.n1 sense_amplifier_0.out1.t1 9.52217
R225 sense_amplifier_0.out1.n1 sense_amplifier_0.out1.t0 9.52217
R226 sense_amplifier_0.out1.n3 sense_amplifier_0.out1 9.08234
R227 sense_amplifier_0.out1 sense_amplifier_0.out1.n8 8.00471
R228 sense_amplifier_0.out1.n8 sense_amplifier_0.out1.n6 4.50239
R229 sense_amplifier_0.out1.n6 sense_amplifier_0.out1.n5 0.898227
R230 sense_amplifier_0.out1.n5 sense_amplifier_0.out1.n4 0.467891
R231 sense_amplifier_0.out1.n4 sense_amplifier_0.out1.n3 0.23963
R232 a_834_510.n2 a_834_510.n1 34.9195
R233 a_834_510.n3 a_834_510.n2 25.5407
R234 a_834_510.n2 a_834_510.n0 25.2907
R235 a_834_510.n1 a_834_510.t1 5.8005
R236 a_834_510.n1 a_834_510.t0 5.8005
R237 a_834_510.n0 a_834_510.t5 5.8005
R238 a_834_510.n0 a_834_510.t4 5.8005
R239 a_834_510.n3 a_834_510.t2 5.8005
R240 a_834_510.t3 a_834_510.n3 5.8005
R241 VDD1.n7 VDD1.n5 1656.75
R242 VDD1.n5 VDD1.n4 1600.08
R243 VDD1.n8 VDD1.t6 196.429
R244 VDD1.n10 VDD1.n4 186.093
R245 VDD1.n6 VDD1.t0 183.929
R246 VDD1.n10 VDD1.n0 176.72
R247 VDD1.t2 VDD1.n7 146.282
R248 VDD1.t4 VDD1.n4 144.881
R249 VDD1.n1 VDD1.t5 85.2064
R250 VDD1.n3 VDD1.t3 84.7281
R251 VDD1.n2 VDD1.t7 84.7281
R252 VDD1.n1 VDD1.t1 84.7281
R253 VDD1.t0 VDD1.t4 78.5719
R254 VDD1.t6 VDD1.t2 78.5719
R255 VDD1.n9 VDD1.n8 38.0519
R256 VDD1.n7 VDD1.n0 16.8187
R257 VDD1.n8 VDD1.n6 12.5005
R258 VDD1.n6 VDD1.n5 6.60764
R259 VDD1.n9 VDD1.n5 5.77063
R260 VDD1.n12 VDD1.n0 1.92668
R261 VDD1.n2 VDD1.n1 0.957022
R262 VDD1.n10 VDD1.n9 0.713588
R263 VDD1.n11 VDD1.n10 0.647749
R264 VDD1.n3 VDD1.n2 0.478761
R265 VDD1 VDD1.n12 0.394487
R266 VDD1.n11 VDD1.n3 0.337457
R267 VDD1.n12 VDD1.n11 0.0804051
R268 nd.n0 nd.t3 784.053
R269 nd.n0 nd.t1 784.053
R270 nd.n1 nd.t0 784.053
R271 nd.n1 nd.t2 784.053
R272 nd.n2 nd.n0 168.659
R273 nd.n2 nd.n1 167.992
R274 nd nd.n2 17.1141
R275 VDD2.n13 VDD2.n7 2143.14
R276 VDD2.n9 VDD2.n8 2138.43
R277 VDD2.n10 VDD2.n8 1486.67
R278 VDD2.n15 VDD2.n6 228.601
R279 VDD2.n14 VDD2.n0 228.1
R280 VDD2.t3 VDD2.n7 169.983
R281 VDD2.t10 VDD2.n9 164.046
R282 VDD2.n14 VDD2.n2 158.578
R283 VDD2.n11 VDD2.t0 143.49
R284 VDD2.n12 VDD2.t7 141.511
R285 VDD2.t12 VDD2.t3 87.0838
R286 VDD2.t2 VDD2.t12 87.0838
R287 VDD2.t7 VDD2.t2 87.0838
R288 VDD2.t0 VDD2.t9 87.0838
R289 VDD2.t9 VDD2.t5 87.0838
R290 VDD2.t5 VDD2.t10 87.0838
R291 VDD2.n18 VDD2.t1 85.0216
R292 VDD2.n3 VDD2.t8 85.0216
R293 VDD2.n19 VDD2.n1 75.5
R294 VDD2.n5 VDD2.n4 75.5
R295 VDD2.n9 VDD2.n0 20.5561
R296 VDD2.n10 VDD2.n2 20.5561
R297 VDD2.n11 VDD2.n10 20.5561
R298 VDD2.n7 VDD2.n6 20.5561
R299 VDD2.n1 VDD2.t6 9.52217
R300 VDD2.n1 VDD2.t11 9.52217
R301 VDD2.n4 VDD2.t4 9.52217
R302 VDD2.n4 VDD2.t13 9.52217
R303 VDD2.n15 VDD2.n13 5.44168
R304 VDD2.n13 VDD2.n12 5.44168
R305 VDD2.n6 VDD2.n5 2.56343
R306 VDD2.n13 VDD2.n8 2.35344
R307 VDD2.n20 VDD2.n0 2.32446
R308 VDD2.n17 VDD2.n2 2.32446
R309 VDD2.n12 VDD2.n11 1.97967
R310 VDD2.n16 VDD2.n15 0.58175
R311 VDD2.n5 VDD2.n3 0.324029
R312 VDD2.n19 VDD2.n18 0.324029
R313 VDD2.n15 VDD2.n14 0.25148
R314 VDD2.n20 VDD2.n19 0.232118
R315 VDD2.n18 VDD2.n17 0.124275
R316 VDD2.n16 VDD2.n3 0.121824
R317 VDD2 VDD2.n20 0.113245
R318 VDD2.n17 VDD2.n16 0.00295098
C0 a_690_n1522# a_958_n952# 0.030392f
C1 sense_amplifier_0.out2 a_1336_n1386# 0.012202f
C2 sense_amplifier_0.out2 nd 0.440678f
C3 a_1336_n952# a_1336_n1386# 0.003413f
C4 clk nd 0.496564f
C5 d a_958_n952# 1.47e-19
C6 VDD2 sense_amplifier_0.out1 1.20128f
C7 sense_amplifier_0.out2 q 0.105071f
C8 clk q 7.9e-20
C9 nq sense_amplifier_0.out1 0.132388f
C10 a_1336_n952# q 0.013457f
C11 a_690_n1522# VDD2 1.43261f
C12 a_1336_n1386# a_1374_n306# 1.02e-19
C13 a_1374_n306# nd 5.04e-20
C14 a_690_n1522# nq 0.014786f
C15 d VDD2 0.006025f
C16 a_658_510# sense_amplifier_0.out1 1.06381f
C17 d nq 0.001059f
C18 a_690_n1522# a_658_510# 2.08e-21
C19 a_1374_n306# q 0.014789f
C20 q a_958_n952# 0.492009f
C21 a_958_n1386# a_958_n952# 0.003413f
C22 d a_658_510# 0.192064f
C23 clk sense_amplifier_0.out2 0.377965f
C24 a_1336_n1386# VDD2 6.18e-19
C25 a_1336_n952# sense_amplifier_0.out2 0.033952f
C26 VDD2 nd 0.010913f
C27 a_1336_n952# clk 9.87e-20
C28 a_690_n1522# sense_amplifier_0.out1 0.196687f
C29 VDD1 sense_amplifier_0.out1 1.36544f
C30 a_1336_n1386# nq 0.174293f
C31 nq nd 1.23e-19
C32 d sense_amplifier_0.out1 0.500493f
C33 q VDD2 0.589355f
C34 a_958_n1386# VDD2 6.18e-19
C35 a_658_510# nd 0.007929f
C36 sense_amplifier_0.out2 a_1374_n306# 0.197072f
C37 sense_amplifier_0.out2 a_958_n952# 0.003664f
C38 a_690_n1522# d 3.84e-19
C39 nq q 0.227882f
C40 d VDD1 0.380532f
C41 clk a_1374_n306# 0.001226f
C42 nq a_958_n1386# 0.005553f
C43 a_1336_n952# a_1374_n306# 0.030083f
C44 nd sense_amplifier_0.out1 0.199846f
C45 a_690_n1522# nd 4.55e-19
C46 VDD1 nd 0.156169f
C47 sense_amplifier_0.out2 VDD2 1.22237f
C48 clk VDD2 0.004202f
C49 q sense_amplifier_0.out1 0.200954f
C50 a_1336_n952# VDD2 0.497547f
C51 a_958_n1386# sense_amplifier_0.out1 0.010872f
C52 sense_amplifier_0.out2 nq 0.231514f
C53 d nd 0.23702f
C54 clk nq 6.62e-20
C55 a_1336_n952# nq 0.504416f
C56 a_690_n1522# q 0.098152f
C57 a_690_n1522# a_958_n1386# 1.02e-19
C58 sense_amplifier_0.out2 a_658_510# 0.09966f
C59 d q 1.13e-20
C60 clk a_658_510# 3.98e-19
C61 a_1374_n306# VDD2 1.41226f
C62 VDD2 a_958_n952# 0.497771f
C63 a_1374_n306# nq 0.100257f
C64 nq a_958_n952# 0.013457f
C65 sense_amplifier_0.out2 sense_amplifier_0.out1 4.28602f
C66 clk sense_amplifier_0.out1 0.140227f
C67 a_1336_n952# sense_amplifier_0.out1 0.003607f
C68 a_1336_n1386# q 0.005553f
C69 a_690_n1522# sense_amplifier_0.out2 0.164202f
C70 sense_amplifier_0.out2 VDD1 1.21676f
C71 q nd 3.6e-19
C72 clk VDD1 2.6112f
C73 sense_amplifier_0.out2 d 0.125784f
C74 clk d 0.119616f
C75 nq VDD2 0.712378f
C76 a_1374_n306# sense_amplifier_0.out1 0.162437f
C77 q a_958_n1386# 0.188081f
C78 a_958_n952# sense_amplifier_0.out1 0.035356f
C79 a_690_n1522# a_1374_n306# 0.005826f
C80 q VSS2 0.725619f
C81 nq VSS2 0.591677f
C82 nd VSS2 2.40742f
C83 d VSS2 2.1265f
C84 clk VSS2 2.935104f
C85 VDD2 VSS2 5.67921f
C86 VDD1 VSS2 4.595867f
C87 a_1336_n1386# VSS2 0.192064f
C88 a_958_n1386# VSS2 0.190559f
C89 a_1336_n952# VSS2 0.023462f
C90 a_958_n952# VSS2 0.024712f
C91 a_1374_n306# VSS2 0.825208f
C92 a_690_n1522# VSS2 0.830819f
C93 a_658_510# VSS2 0.354057f
C94 sense_amplifier_0.out1 VSS2 5.579126f
C95 sense_amplifier_0.out2 VSS2 5.966842f
C96 VDD1.n0 VSS2 0.04434f
C97 VDD1.t3 VSS2 0.032405f
C98 VDD1.t7 VSS2 0.032405f
C99 VDD1.t1 VSS2 0.032405f
C100 VDD1.t5 VSS2 0.032725f
C101 VDD1.n1 VSS2 0.120595f
C102 VDD1.n2 VSS2 0.063955f
C103 VDD1.n3 VSS2 0.059795f
C104 VDD1.n4 VSS2 0.20253f
C105 VDD1.n5 VSS2 0.182324f
C106 VDD1.t4 VSS2 0.140567f
C107 VDD1.t0 VSS2 0.155433f
C108 VDD1.n6 VSS2 0.116311f
C109 VDD1.n7 VSS2 0.148519f
C110 VDD1.t2 VSS2 0.138805f
C111 VDD1.t6 VSS2 0.162835f
C112 VDD1.n8 VSS2 0.318725f
C113 VDD1.n9 VSS2 0.030449f
C114 VDD1.n10 VSS2 0.306628f
C115 VDD1.n11 VSS2 0.169656f
C116 VDD1.n12 VSS2 0.069497f
C117 a_834_510.t2 VSS2 0.059028f
C118 a_834_510.t5 VSS2 0.059028f
C119 a_834_510.t4 VSS2 0.059028f
C120 a_834_510.n0 VSS2 0.136068f
C121 a_834_510.t1 VSS2 0.059028f
C122 a_834_510.t0 VSS2 0.059028f
C123 a_834_510.n1 VSS2 0.258102f
C124 a_834_510.n2 VSS2 1.11221f
C125 a_834_510.n3 VSS2 0.139449f
C126 a_834_510.t3 VSS2 0.059028f
C127 sense_amplifier_0.out1.t10 VSS2 0.059931f
C128 sense_amplifier_0.out1.t7 VSS2 0.025764f
C129 sense_amplifier_0.out1.n0 VSS2 0.072496f
C130 sense_amplifier_0.out1.t1 VSS2 0.033915f
C131 sense_amplifier_0.out1.t0 VSS2 0.033915f
C132 sense_amplifier_0.out1.n1 VSS2 0.07124f
C133 sense_amplifier_0.out1.t3 VSS2 0.126387f
C134 sense_amplifier_0.out1.t2 VSS2 0.124707f
C135 sense_amplifier_0.out1.t6 VSS2 0.054731f
C136 sense_amplifier_0.out1.t4 VSS2 0.024932f
C137 sense_amplifier_0.out1.n2 VSS2 0.060896f
C138 sense_amplifier_0.out1.n3 VSS2 0.412182f
C139 sense_amplifier_0.out1.n4 VSS2 0.249269f
C140 sense_amplifier_0.out1.n5 VSS2 0.238209f
C141 sense_amplifier_0.out1.t8 VSS2 0.067054f
C142 sense_amplifier_0.out1.n6 VSS2 0.087045f
C143 sense_amplifier_0.out1.t5 VSS2 0.051106f
C144 sense_amplifier_0.out1.t9 VSS2 0.056624f
C145 sense_amplifier_0.out1.n7 VSS2 0.067437f
C146 sense_amplifier_0.out1.n8 VSS2 0.776775f
C147 sense_amplifier_0.out2.n0 VSS2 0.489902f
C148 sense_amplifier_0.out2.n1 VSS2 0.600837f
C149 sense_amplifier_0.out2.t5 VSS2 0.0562f
C150 sense_amplifier_0.out2.t4 VSS2 0.025601f
C151 sense_amplifier_0.out2.n2 VSS2 0.062604f
C152 sense_amplifier_0.out2.t2 VSS2 0.034825f
C153 sense_amplifier_0.out2.t3 VSS2 0.034825f
C154 sense_amplifier_0.out2.n3 VSS2 0.073891f
C155 sense_amplifier_0.out2.t1 VSS2 0.129471f
C156 sense_amplifier_0.out2.t10 VSS2 0.06154f
C157 sense_amplifier_0.out2.t7 VSS2 0.026455f
C158 sense_amplifier_0.out2.n4 VSS2 0.074526f
C159 sense_amplifier_0.out2.t9 VSS2 0.069659f
C160 sense_amplifier_0.out2.t6 VSS2 0.052477f
C161 sense_amplifier_0.out2.t8 VSS2 0.058144f
C162 sense_amplifier_0.out2.n5 VSS2 0.068475f
C163 sense_amplifier_0.out2.t0 VSS2 0.129471f
C164 sense_amplifier_0.out2.n6 VSS2 0.483754f
C165 a_570_510.t4 VSS2 0.024913f
C166 a_570_510.t5 VSS2 0.024913f
C167 a_570_510.t3 VSS2 0.024913f
C168 a_570_510.n0 VSS2 0.060114f
C169 a_570_510.t6 VSS2 0.024913f
C170 a_570_510.t2 VSS2 0.024913f
C171 a_570_510.n1 VSS2 0.060114f
C172 a_570_510.t9 VSS2 0.024913f
C173 a_570_510.t11 VSS2 0.024913f
C174 a_570_510.n2 VSS2 0.057409f
C175 a_570_510.t8 VSS2 0.024913f
C176 a_570_510.t10 VSS2 0.024913f
C177 a_570_510.n3 VSS2 0.060272f
C178 a_570_510.n4 VSS2 0.340434f
C179 a_570_510.t7 VSS2 0.024913f
C180 a_570_510.t12 VSS2 0.024913f
C181 a_570_510.n5 VSS2 0.052659f
C182 a_570_510.n6 VSS2 0.140942f
C183 a_570_510.n7 VSS2 0.22019f
C184 a_570_510.n8 VSS2 0.182473f
C185 a_570_510.t1 VSS2 0.097139f
C186 a_570_510.n9 VSS2 0.369186f
C187 a_570_510.n10 VSS2 0.060114f
C188 a_570_510.t0 VSS2 0.024913f
C189 clk.t3 VSS2 0.074319f
C190 clk.t2 VSS2 0.074152f
C191 clk.n0 VSS2 0.319828f
C192 clk.t0 VSS2 0.057095f
C193 clk.t4 VSS2 0.057095f
C194 clk.t1 VSS2 0.057095f
C195 clk.t5 VSS2 0.057095f
C196 clk.t6 VSS2 0.06326f
C197 clk.n1 VSS2 0.055633f
C198 clk.n2 VSS2 0.032794f
C199 clk.n3 VSS2 0.032794f
C200 clk.n4 VSS2 0.049399f
C201 clk.n5 VSS2 0.742826f
.ends

