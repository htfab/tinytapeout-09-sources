magic
tech sky130A
magscale 1 2
timestamp 1730183176
<< nwell >>
rect 2916 3096 3084 3616
rect 2916 2868 3076 3096
rect 2916 2648 3084 2868
rect 3396 2648 3456 3616
rect 4320 -190 4498 -116
<< pwell >>
rect 3076 1732 3090 1794
rect 3820 1718 3886 1784
rect 2796 532 2862 598
rect 2420 -1680 2504 -1390
rect 2692 -1514 2760 -1396
rect 2800 -1514 2870 -1492
rect 2692 -1544 3906 -1514
rect 2682 -1552 3906 -1544
rect 3960 -1552 3966 -1514
rect 4216 -1548 4282 -1492
rect 4532 -1548 4598 -1492
rect 2682 -1558 3966 -1552
rect 2682 -1646 2754 -1558
rect 2800 -1930 2870 -1558
rect 4678 -1672 4762 -1382
rect 4848 -1548 4914 -1492
<< poly >>
rect 3742 1642 3964 1708
rect 2622 1442 2844 1508
rect 2604 532 2862 598
rect 3120 532 3378 598
<< locali >>
rect 2404 3780 3776 3818
rect 2404 3648 2430 3780
rect 3748 3648 3776 3780
rect 2404 3580 3776 3648
rect 2910 1648 2988 2596
rect 2458 1594 3578 1648
rect 2604 548 2862 582
rect 3524 446 3578 1594
rect 2420 424 4128 446
rect 2420 264 2452 424
rect 4100 264 4128 424
rect 2420 244 4128 264
rect 2098 138 5094 172
rect 2098 2 2144 138
rect 5052 2 5094 138
rect 2098 -48 5094 2
rect 2100 -1686 5092 -1634
rect 2100 -1800 2120 -1686
rect 5072 -1800 5092 -1686
rect 2100 -1816 5092 -1800
<< viali >>
rect 2430 3648 3748 3780
rect 2452 264 4100 424
rect 2144 2 5052 138
rect 2120 -1800 5072 -1686
<< metal1 >>
rect 2206 3780 3776 3818
rect 2206 3648 2430 3780
rect 3748 3690 3776 3780
rect 3748 3648 5094 3690
rect 2206 3616 5094 3648
rect 2286 3396 2346 3616
rect 2374 3426 2384 3494
rect 2450 3426 2460 3494
rect 3522 3428 3532 3494
rect 3598 3428 3608 3494
rect 3636 3396 3696 3616
rect 2286 3162 2350 3396
rect 3632 3186 3696 3396
rect 2798 3096 3184 3166
rect 2476 2868 2666 3096
rect 2754 3070 3184 3096
rect 3312 3070 3498 3168
rect 2754 2868 2800 3070
rect 2476 2796 2560 2868
rect 2498 2782 2560 2796
rect 2498 2728 2504 2782
rect 2174 2658 2244 2664
rect 2174 2606 2184 2658
rect 2174 662 2244 2606
rect 2498 2500 2560 2728
rect 2174 610 2182 662
rect 2236 610 2244 662
rect 2174 604 2244 610
rect 2288 2432 2560 2500
rect 2700 2658 2766 2828
rect 2700 2604 2708 2658
rect 2700 2454 2766 2604
rect 3216 2782 3282 2828
rect 3274 2728 3282 2782
rect 3216 2454 3282 2728
rect 3312 2658 3374 3070
rect 3368 2604 3374 2658
rect 3312 2498 3374 2604
rect 3474 2546 3480 2608
rect 3532 2546 4914 2608
rect 3474 2540 4914 2546
rect 2288 662 2358 2432
rect 2498 2422 2560 2432
rect 3312 2432 4598 2498
rect 2498 2416 2622 2422
rect 2748 2416 2810 2422
rect 2498 2194 2564 2416
rect 2618 2194 2628 2416
rect 2744 2194 2754 2416
rect 2808 2194 2810 2416
rect 3068 2416 3142 2422
rect 3312 2416 3374 2432
rect 3068 2194 3078 2416
rect 3132 2194 3142 2416
rect 3260 2194 3270 2416
rect 3324 2194 3374 2416
rect 2560 2188 2622 2194
rect 2748 2188 2810 2194
rect 2480 2050 2538 2056
rect 2480 1828 2486 2050
rect 2480 1420 2538 1828
rect 2652 2050 2718 2056
rect 2652 1828 2658 2050
rect 2710 1828 2718 2050
rect 2652 1822 2718 1828
rect 2996 2050 3054 2056
rect 2996 1828 3002 2050
rect 2604 1734 2670 1790
rect 2700 1502 2766 1508
rect 2700 1450 2706 1502
rect 2760 1450 2766 1502
rect 2700 1448 2766 1450
rect 2996 1420 3054 1828
rect 3168 2050 3234 2058
rect 3168 1828 3174 2050
rect 3226 1828 3234 2050
rect 3168 1822 3234 1828
rect 3120 1734 3186 1790
rect 3820 1652 3826 1708
rect 3880 1652 3886 1708
rect 3774 1614 3836 1620
rect 3216 1452 3282 1508
rect 2480 1414 2620 1420
rect 2480 1192 2562 1414
rect 2616 1192 2620 1414
rect 2480 1186 2620 1192
rect 2750 1414 2812 1420
rect 2750 1192 2754 1414
rect 2808 1192 2812 1414
rect 2750 1186 2812 1192
rect 2996 1414 3136 1420
rect 2996 1192 3078 1414
rect 3132 1192 3136 1414
rect 2996 1186 3136 1192
rect 3266 1414 3328 1420
rect 3266 1192 3270 1414
rect 3324 1192 3328 1414
rect 3774 1392 3778 1614
rect 3832 1392 3836 1614
rect 3774 1386 3836 1392
rect 3966 1614 4028 1620
rect 3966 1392 3970 1614
rect 4024 1392 4028 1614
rect 3966 1386 4028 1392
rect 3266 1186 3328 1192
rect 2288 610 2296 662
rect 2350 610 2358 662
rect 2654 848 2716 854
rect 2654 626 2658 848
rect 2712 626 2716 848
rect 2654 620 2716 626
rect 2846 848 2908 854
rect 2846 626 2850 848
rect 2904 626 2908 848
rect 2846 620 2908 626
rect 3170 848 3232 854
rect 3170 626 3174 848
rect 3228 626 3232 848
rect 3170 620 3232 626
rect 3362 848 3424 854
rect 3362 626 3366 848
rect 3420 626 3424 848
rect 3362 620 3424 626
rect 3678 848 3740 854
rect 3678 626 3682 848
rect 3736 626 3740 848
rect 3678 620 3740 626
rect 3870 848 3932 854
rect 3870 626 3874 848
rect 3928 626 3932 848
rect 3870 620 3932 626
rect 2288 604 2358 610
rect 2604 542 2862 588
rect 3120 536 3128 588
rect 3370 536 3378 588
rect 3120 532 3378 536
rect 3724 532 3790 588
rect 3916 532 3982 588
rect 4020 446 4074 774
rect 4532 668 4598 2432
rect 4532 614 4538 668
rect 4592 614 4598 668
rect 4532 608 4598 614
rect 4848 666 4914 2540
rect 4848 614 4854 666
rect 4908 614 4914 666
rect 4848 608 4914 614
rect 2156 444 4128 446
rect 1956 424 4128 444
rect 1956 264 2452 424
rect 4100 264 4128 424
rect 1956 244 4128 264
rect 2014 -1670 2068 244
rect 5010 172 5094 3616
rect 2100 138 5094 172
rect 2100 2 2144 138
rect 5052 2 5094 138
rect 2100 -14 5094 2
rect 2276 -134 2342 -130
rect 2276 -186 2282 -134
rect 2336 -186 2342 -134
rect 2276 -190 2342 -186
rect 2376 -490 2430 -14
rect 3224 -124 3304 -116
rect 2592 -136 2658 -134
rect 2592 -188 2598 -136
rect 2652 -188 2658 -136
rect 2592 -190 2658 -188
rect 2908 -190 2974 -134
rect 3224 -182 3232 -124
rect 3296 -182 3304 -124
rect 3224 -190 3304 -182
rect 2376 -560 2562 -490
rect 2692 -560 2878 -490
rect 3006 -560 3192 -490
rect 3566 -498 3620 -14
rect 4320 -124 4498 -116
rect 3900 -190 3966 -134
rect 4216 -190 4282 -134
rect 4320 -182 4330 -124
rect 4392 -182 4498 -124
rect 4320 -190 4498 -182
rect 4532 -122 4598 -116
rect 4532 -184 4538 -122
rect 4592 -184 4598 -122
rect 4532 -190 4598 -184
rect 4436 -360 4498 -190
rect 3320 -562 3870 -498
rect 4760 -512 4814 -14
rect 4848 -122 4914 -116
rect 4848 -184 4854 -122
rect 4908 -184 4914 -122
rect 4848 -190 4914 -184
rect 3994 -582 4188 -512
rect 4310 -582 4504 -512
rect 4626 -582 4820 -512
rect 2182 -1116 2242 -642
rect 2182 -1170 2188 -1116
rect 2182 -1460 2242 -1170
rect 2276 -1228 2342 -872
rect 2592 -1020 2658 -870
rect 2592 -1072 2600 -1020
rect 2592 -1078 2658 -1072
rect 2592 -1164 2658 -1158
rect 2592 -1222 2598 -1164
rect 2652 -1222 2658 -1164
rect 2592 -1228 2658 -1222
rect 2692 -1326 2744 -720
rect 2908 -878 2974 -872
rect 2908 -932 2914 -878
rect 2968 -932 2974 -878
rect 2908 -938 2974 -932
rect 2802 -1020 2974 -1014
rect 2858 -1072 2974 -1020
rect 2802 -1078 2974 -1072
rect 2908 -1228 2974 -1078
rect 3224 -1228 3290 -872
rect 3900 -1228 3966 -872
rect 4216 -878 4282 -872
rect 4216 -930 4222 -878
rect 4276 -930 4282 -878
rect 4216 -936 4282 -930
rect 4216 -1022 4402 -1016
rect 4216 -1074 4342 -1022
rect 4396 -1074 4402 -1022
rect 4216 -1080 4402 -1074
rect 4216 -1228 4282 -1080
rect 4440 -1322 4498 -718
rect 4532 -1022 4598 -872
rect 4532 -1074 4538 -1022
rect 4592 -1074 4598 -1022
rect 4532 -1080 4598 -1074
rect 4532 -1170 4598 -1164
rect 4532 -1222 4538 -1170
rect 4592 -1222 4598 -1170
rect 4532 -1228 4598 -1222
rect 4848 -1228 4914 -872
rect 4948 -1112 5006 -680
rect 4948 -1120 5020 -1112
rect 4948 -1176 4956 -1120
rect 5012 -1176 5020 -1120
rect 4948 -1184 5020 -1176
rect 2372 -1396 2558 -1326
rect 2692 -1396 2878 -1326
rect 2276 -1548 2342 -1492
rect 2420 -1670 2504 -1396
rect 2592 -1548 2658 -1492
rect 2692 -1498 2760 -1396
rect 3006 -1398 3192 -1328
rect 3320 -1398 3870 -1334
rect 3994 -1392 4188 -1322
rect 4310 -1330 4504 -1322
rect 4310 -1386 4434 -1330
rect 4488 -1386 4504 -1330
rect 4310 -1392 4504 -1386
rect 4626 -1392 4820 -1322
rect 4948 -1380 5006 -1184
rect 2692 -1552 2698 -1498
rect 2908 -1548 2974 -1492
rect 3224 -1548 3290 -1492
rect 2692 -1558 2760 -1552
rect 3550 -1670 3634 -1398
rect 3900 -1498 3966 -1492
rect 3900 -1554 3906 -1498
rect 3960 -1554 3966 -1498
rect 4216 -1548 4282 -1492
rect 4532 -1548 4598 -1492
rect 3900 -1558 3966 -1554
rect 4678 -1670 4762 -1392
rect 4848 -1548 4914 -1492
rect 2014 -1686 5092 -1670
rect 2014 -1800 2120 -1686
rect 5072 -1800 5092 -1686
rect 2014 -1816 5092 -1800
<< via1 >>
rect 2384 3426 2450 3494
rect 3532 3428 3598 3494
rect 2504 2728 2560 2782
rect 2184 2606 2244 2658
rect 2182 610 2236 662
rect 2708 2604 2766 2658
rect 3216 2728 3274 2782
rect 3312 2604 3368 2658
rect 3480 2546 3532 2608
rect 2564 2194 2618 2416
rect 2754 2194 2808 2416
rect 3078 2194 3132 2416
rect 3270 2194 3324 2416
rect 2486 1828 2538 2050
rect 2658 1828 2710 2050
rect 3002 1828 3054 2050
rect 2706 1450 2760 1502
rect 3174 1828 3226 2050
rect 3826 1652 3880 1708
rect 2562 1192 2616 1414
rect 2754 1192 2808 1414
rect 3078 1192 3132 1414
rect 3270 1192 3324 1414
rect 3778 1392 3832 1614
rect 3970 1392 4024 1614
rect 2296 610 2350 662
rect 2658 626 2712 848
rect 2850 626 2904 848
rect 3174 626 3228 848
rect 3366 626 3420 848
rect 3682 626 3736 848
rect 3874 626 3928 848
rect 3128 536 3370 588
rect 4538 614 4592 668
rect 4854 614 4908 666
rect 2282 -186 2336 -134
rect 2598 -188 2652 -136
rect 3232 -182 3296 -124
rect 4330 -182 4392 -124
rect 4538 -184 4592 -122
rect 4854 -184 4908 -122
rect 2188 -1170 2242 -1116
rect 2600 -1072 2658 -1020
rect 2598 -1222 2652 -1164
rect 2914 -932 2968 -878
rect 2802 -1072 2858 -1020
rect 4222 -930 4276 -878
rect 4342 -1074 4396 -1022
rect 4538 -1074 4592 -1022
rect 4538 -1222 4592 -1170
rect 4956 -1176 5012 -1120
rect 4434 -1386 4488 -1330
rect 2698 -1552 2760 -1498
rect 3906 -1554 3960 -1498
<< metal2 >>
rect 2060 3930 2260 4130
rect 2384 3930 2584 4130
rect 2060 1508 2132 3930
rect 2384 3504 2450 3930
rect 4182 3928 4382 4128
rect 2384 3494 3886 3504
rect 2450 3428 3532 3494
rect 3598 3428 3886 3494
rect 2450 3426 3886 3428
rect 2384 3418 3886 3426
rect 2384 3416 2450 3418
rect 2498 2782 3536 2786
rect 2498 2728 2504 2782
rect 2560 2728 3216 2782
rect 3274 2728 3536 2782
rect 2498 2724 3536 2728
rect 2174 2658 3374 2664
rect 2174 2606 2184 2658
rect 2244 2606 2708 2658
rect 2174 2604 2708 2606
rect 2766 2604 3312 2658
rect 3368 2604 3374 2658
rect 2174 2600 3374 2604
rect 3474 2608 3536 2724
rect 3474 2546 3480 2608
rect 3532 2546 3536 2608
rect 3474 2540 3536 2546
rect 2564 2422 2618 2426
rect 2754 2422 2808 2426
rect 2560 2416 2810 2422
rect 2560 2194 2564 2416
rect 2618 2194 2754 2416
rect 2808 2194 2810 2416
rect 2560 2188 2810 2194
rect 3078 2416 3132 2426
rect 3270 2416 3324 2426
rect 3132 2194 3270 2416
rect 2564 2184 2618 2188
rect 2754 2184 2808 2188
rect 3078 2184 3132 2194
rect 3270 2184 3324 2194
rect 2480 2050 2718 2056
rect 2480 1828 2486 2050
rect 2538 1828 2658 2050
rect 2710 1828 2718 2050
rect 2480 1822 2718 1828
rect 2996 2050 3234 2056
rect 2996 1828 3002 2050
rect 3054 1828 3174 2050
rect 3226 1828 3234 2050
rect 2996 1822 3234 1828
rect 3820 1708 3886 3418
rect 3820 1652 3826 1708
rect 3880 1652 3886 1708
rect 3774 1614 4028 1620
rect 2060 1502 2766 1508
rect 2060 1450 2706 1502
rect 2760 1450 2766 1502
rect 2060 1448 2766 1450
rect 2558 1414 2812 1420
rect 2558 1192 2562 1414
rect 2616 1192 2754 1414
rect 2808 1192 2812 1414
rect 2558 1186 2812 1192
rect 3074 1414 3328 1420
rect 3074 1192 3078 1414
rect 3132 1192 3270 1414
rect 3324 1192 3328 1414
rect 3774 1392 3778 1614
rect 3832 1392 3970 1614
rect 4024 1392 4028 1614
rect 3774 1386 4028 1392
rect 3074 1186 3328 1192
rect 2654 848 3932 854
rect 2174 662 2246 670
rect 2174 610 2182 662
rect 2236 610 2246 662
rect 2174 -130 2246 610
rect 2288 662 2358 670
rect 2288 610 2296 662
rect 2350 610 2358 662
rect 2654 626 2658 848
rect 2712 626 2850 848
rect 2904 626 3174 848
rect 3228 626 3366 848
rect 3420 626 3682 848
rect 3736 626 3874 848
rect 3928 626 3932 848
rect 2654 620 3932 626
rect 2288 124 2358 610
rect 3120 536 3128 588
rect 3370 536 3378 588
rect 3120 532 3378 536
rect 4182 532 4250 3928
rect 3120 480 4250 532
rect 4532 668 4598 674
rect 4532 614 4538 668
rect 4592 614 4598 668
rect 2288 54 2658 124
rect 2174 -134 2342 -130
rect 2174 -186 2282 -134
rect 2336 -186 2342 -134
rect 2174 -190 2342 -186
rect 2592 -136 2658 54
rect 2592 -188 2598 -136
rect 2652 -188 2658 -136
rect 2592 -190 2658 -188
rect 3224 -124 4400 -116
rect 3224 -182 3232 -124
rect 3296 -182 4330 -124
rect 4392 -182 4400 -124
rect 3224 -190 4400 -182
rect 4532 -122 4598 614
rect 4532 -184 4538 -122
rect 4592 -184 4598 -122
rect 4532 -190 4598 -184
rect 4848 666 4914 672
rect 4848 614 4854 666
rect 4908 614 4914 666
rect 4848 -122 4914 614
rect 4848 -184 4854 -122
rect 4908 -184 4914 -122
rect 4848 -190 4914 -184
rect 2908 -878 3040 -872
rect 2908 -932 2914 -878
rect 2968 -932 3040 -878
rect 2908 -938 3040 -932
rect 2592 -1020 2862 -1014
rect 2592 -1072 2600 -1020
rect 2658 -1072 2802 -1020
rect 2858 -1072 2862 -1020
rect 2592 -1078 2862 -1072
rect 2974 -1110 3040 -938
rect 2182 -1116 3040 -1110
rect 2182 -1170 2188 -1116
rect 2242 -1164 3040 -1116
rect 2242 -1170 2598 -1164
rect 2182 -1176 2598 -1170
rect 2592 -1222 2598 -1176
rect 2652 -1176 3040 -1164
rect 4152 -878 4282 -872
rect 4152 -930 4222 -878
rect 4276 -930 4282 -878
rect 4152 -936 4282 -930
rect 4152 -1112 4216 -936
rect 4336 -1022 4598 -1016
rect 4336 -1074 4342 -1022
rect 4396 -1074 4538 -1022
rect 4592 -1074 4598 -1022
rect 4336 -1080 4598 -1074
rect 4152 -1120 5020 -1112
rect 4152 -1170 4956 -1120
rect 4152 -1172 4538 -1170
rect 2652 -1222 2658 -1176
rect 2592 -1228 2658 -1222
rect 4532 -1222 4538 -1172
rect 4592 -1172 4956 -1170
rect 4592 -1222 4598 -1172
rect 4948 -1176 4956 -1172
rect 5012 -1176 5020 -1120
rect 4948 -1184 5020 -1176
rect 4532 -1228 4598 -1222
rect 4428 -1330 4498 -1322
rect 4428 -1386 4434 -1330
rect 4488 -1386 4498 -1330
rect 2692 -1498 3966 -1492
rect 2692 -1552 2698 -1498
rect 2760 -1552 3906 -1498
rect 2692 -1554 3906 -1552
rect 3960 -1554 3966 -1498
rect 2692 -1558 3966 -1554
rect 2800 -1930 2870 -1558
rect 2670 -2130 2870 -1930
rect 4428 -1922 4498 -1386
rect 4428 -2122 4628 -1922
use sky130_fd_pr__nfet_01v8_95PS5T  sky130_fd_pr__nfet_01v8_95PS5T_0
timestamp 1730034632
transform 1 0 2733 0 1 1020
box -311 -610 311 610
use sky130_fd_pr__nfet_01v8_648S5X  sky130_fd_pr__nfet_01v8_648S5X_0
timestamp 1730034632
transform 1 0 2309 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_LGES5M  sky130_fd_pr__nfet_01v8_LGES5M_0
timestamp 1730034632
transform 1 0 2685 0 1 2122
box -263 -510 263 510
use sky130_fd_pr__pfet_01v8_MGSNAN  sky130_fd_pr__pfet_01v8_MGSNAN_0
timestamp 1730064633
transform 1 0 2417 0 1 3132
box -211 -484 211 484
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1730034632
transform 1 0 3933 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_MGSNAN  XM4
timestamp 1730064633
transform 1 0 3565 0 1 3132
box -211 -484 211 484
use sky130_fd_pr__pfet_01v8_LGSNAL  XM5
timestamp 1730064633
transform 1 0 3249 0 1 3132
box -211 -484 211 484
use sky130_fd_pr__pfet_01v8_LGSNAL  XM6
timestamp 1730064633
transform 1 0 2733 0 1 3132
box -211 -484 211 484
use sky130_fd_pr__nfet_01v8_LGES5M  XM7
timestamp 1730034632
transform 1 0 3201 0 1 2122
box -263 -510 263 510
use sky130_fd_pr__nfet_01v8_84PS53  XM9
timestamp 1730034632
transform 1 0 3853 0 1 1120
box -311 -710 311 710
use sky130_fd_pr__nfet_01v8_95PS5T  XM10
timestamp 1730034632
transform 1 0 3249 0 1 1020
box -311 -610 311 610
use sky130_fd_pr__pfet_01v8_XGSNAL  XM12
timestamp 1730034632
transform 1 0 4881 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM13
timestamp 1730034632
transform 1 0 4881 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XM14
timestamp 1730034632
transform 1 0 2309 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM16
timestamp 1730034632
transform 1 0 2625 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM17
timestamp 1730034632
transform 1 0 2625 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XM18
timestamp 1730034632
transform 1 0 4565 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM19
timestamp 1730034632
transform 1 0 4565 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XM20
timestamp 1730034632
transform 1 0 3933 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM21
timestamp 1730034632
transform 1 0 4249 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM22
timestamp 1730034632
transform 1 0 2941 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XGSNAL  XM23
timestamp 1730034632
transform 1 0 3257 0 1 -531
box -211 -519 211 519
use sky130_fd_pr__nfet_01v8_648S5X  XM24
timestamp 1730034632
transform 1 0 2941 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM25
timestamp 1730034632
transform 1 0 4249 0 1 -1360
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM26
timestamp 1730034632
transform 1 0 3257 0 1 -1360
box -211 -310 211 310
<< labels >>
flabel metal1 2206 3618 2406 3818 0 FreeSans 256 0 0 0 VDD
port 5 nsew
flabel metal1 1956 244 2156 444 0 FreeSans 256 0 0 0 VSS
port 6 nsew
flabel metal2 2060 3930 2260 4130 0 FreeSans 256 0 0 0 d
port 0 nsew
flabel metal2 2384 3930 2584 4130 0 FreeSans 256 0 0 0 clk
port 2 nsew
flabel metal2 4182 3928 4382 4128 0 FreeSans 256 0 0 0 nd
port 1 nsew
flabel metal2 2670 -2130 2870 -1930 0 FreeSans 256 0 0 0 q
port 3 nsew
flabel metal2 4428 -2122 4628 -1922 0 FreeSans 256 0 0 0 nq
port 4 nsew
<< end >>
