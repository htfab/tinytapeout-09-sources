* NGSPICE file created from tdc_parax.ext - technology: sky130A

.subckt tdc_parax term_4 stop term_3 term_5 term_2 term_1 term_6 term_0 term_7 start
+ VSS VDD
X0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VDD.t365 VDD.t364 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1 a_17444_296# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 term_7.t3 VSS.t380 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X2 a_14862_2192# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 a_14774_2192.t10 VSS.t382 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X3 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8732_1376# a_8694_730# VDD.t224 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X4 diff_gen_0.delay_unit_2_6.in_1.t2 diff_gen_0.delay_unit_2_5.in_2.t8 VSS.t437 VSS.t436 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X5 VDD.t503 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDD.t502 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 a_4130_296# VSS.t581 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X7 a_12492_2192.t9 vernier_delay_line_0.stop_strong.t32 VSS.t135 VSS.t134 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X8 VSS.t563 diff_gen_0.delay_unit_2_2.in_1.t8 diff_gen_0.delay_unit_2_3.in_2.t2 VSS.t562 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X9 VDD.t31 start_buffer_0.start_buff.t10 start_buffer_0.start_delay.t7 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 VSS.t457 VSS.t456 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X11 a_n6458_3464.t3 a_n6748_3464# VSS.t234 VSS.t233 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 VSS.t92 diff_gen_0.delay_unit_2_1.in_2.t8 diff_gen_0.delay_unit_2_1.in_1.t0 VSS.t91 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X13 VSS.t69 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 VSS.t68 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X14 diff_gen_0.delay_unit_2_5.in_2.t7 diff_gen_0.delay_unit_2_4.in_1.t8 VSS.t550 VSS.t549 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X15 vernier_delay_line_0.start_neg.t2 diff_gen_0.delay_unit_2_6.in_1.t8 VSS.t156 VSS.t155 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X16 a_5910_2192.t5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 a_5646_2192.t9 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X17 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X18 a_13258_296# term_5.t4 VSS.t148 VSS.t147 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X19 start_buffer_0.start_buff.t3 a_n11872_5654# VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X20 a_3364_2192.t10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 a_3452_2192# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X21 VDD.t134 diff_gen_0.delay_unit_2_5.in_2.t9 diff_gen_0.delay_unit_2_5.in_1.t4 VDD.t133 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X22 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 a_1848_296# VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X23 a_3364_2192.t6 vernier_delay_line_0.stop_strong.t33 VSS.t133 VSS.t132 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X24 a_14774_2192.t6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 a_15038_2192.t5 VSS.t334 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X25 VSS.t353 vernier_delay_line_0.stop_strong.t34 a_1082_2192.t8 VSS.t352 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X26 VSS.t88 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 VSS.t87 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X27 vernier_delay_line_0.delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X28 VDD.t339 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VDD.t338 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X29 VDD.t388 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8316_730# VDD.t387 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X30 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 VSS.t336 VSS.t335 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X31 a_14774_2192.t11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 a_15038_2192.t4 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X32 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VDD.t416 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X33 VDD.t45 diff_gen_0.delay_unit_2_3.in_2.t8 diff_gen_0.delay_unit_2_4.in_1.t6 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X34 VSS.t542 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VSS.t541 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X35 a_15578_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VSS.t388 VSS.t387 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X36 VDD.t472 diff_gen_0.delay_unit_2_5.in_1.t8 diff_gen_0.delay_unit_2_6.in_2.t7 VDD.t471 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X37 diff_gen_0.delay_unit_2_1.in_2.t6 start_buffer_0.start_buff.t11 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X38 VDD.t414 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X39 a_8016_2192# vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 a_7928_2192.t3 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X40 a_17444_730# a_17176_160# term_7.t0 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X41 VDD.t295 vernier_delay_line_0.start_pos.t8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X42 diff_gen_0.delay_unit_2_1.in_1.t7 start_buffer_0.start_delay.t8 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X43 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VSS.t150 VSS.t149 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X44 VDD.t437 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X45 a_5646_2192.t4 vernier_delay_line_0.stop_strong.t35 VSS.t348 VSS.t347 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X46 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_4168_1376# a_4130_730# VDD.t494 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X47 VSS.t261 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1470_296# VSS.t260 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X48 VSS.t342 vernier_delay_line_0.stop_strong.t36 a_3364_2192.t5 VSS.t341 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X49 VDD.t317 diff_gen_0.delay_unit_2_2.in_2.t8 diff_gen_0.delay_unit_2_3.in_1.t5 VDD.t316 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X50 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 VSS.t355 VSS.t354 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X51 VSS.t346 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 a_12612_160# VSS.t345 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X52 VDD.t451 vernier_delay_line_0.start_neg.t8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 VDD.t450 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X53 a_17056_2192.t3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 a_17144_2192# VSS.t440 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X54 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 vernier_delay_line_0.stop_strong.t37 VDD.t313 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X55 VDD.t101 diff_gen_0.delay_unit_2_3.in_1.t8 diff_gen_0.delay_unit_2_3.in_2.t7 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X56 a_17056_2192.t12 vernier_delay_line_0.stop_strong.t38 VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X57 vernier_delay_line_0.start_pos.t4 diff_gen_0.delay_unit_2_6.in_2.t8 VSS.t427 VSS.t426 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X58 VSS.t279 a_6450_1376# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VSS.t278 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X59 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 VSS.t190 VSS.t189 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X60 VDD.t12 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X61 a_13258_730# term_5.t5 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X62 a_10210_2192.t3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 a_10474_2192.t2 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X63 a_1170_2192# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X64 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1886_1376# a_1848_730# VDD.t180 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X65 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 VDD.t325 VDD.t324 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X66 a_7928_2192.t12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 a_8192_2192.t5 VSS.t488 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X67 VDD.t259 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 VDD.t258 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X68 a_12756_2192.t5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X69 VSS.t485 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15162_296# VSS.t484 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X70 a_1082_2192.t12 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 a_1170_2192# VSS.t531 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X71 a_15578_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VDD.t363 VDD.t362 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X72 a_7928_2192.t9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 a_8192_2192.t4 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X73 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X74 VDD.t63 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X75 VSS.t176 diff_gen_0.delay_unit_2_1.in_1.t8 diff_gen_0.delay_unit_2_2.in_2.t4 VSS.t175 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X76 a_1082_2192.t7 vernier_delay_line_0.stop_strong.t39 VSS.t338 VSS.t337 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X77 VDD.t165 vernier_delay_line_0.stop_strong.t40 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X78 VSS.t90 start_buffer_0.start_delay.t9 start_buffer_0.start_buff.t8 VSS.t89 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X79 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 VSS.t570 VSS.t569 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X80 VDD.t253 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 VDD.t252 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X81 a_12492_2192.t0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 a_12580_2192# VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X82 a_n6458_3464.t7 a_n6748_3464# VDD.t205 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X83 VSS.t291 diff_gen_0.delay_unit_2_1.in_2.t9 diff_gen_0.delay_unit_2_2.in_1.t5 VSS.t290 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X84 VDD.t234 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1470_730# VDD.t233 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X85 VSS.t188 vernier_delay_line_0.stop_strong.t41 a_10210_2192.t12 VSS.t187 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X86 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 a_10976_296# VSS.t468 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X87 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VSS.t312 VSS.t311 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X88 VDD.t466 diff_gen_0.delay_unit_2_4.in_2.t8 diff_gen_0.delay_unit_2_4.in_1.t7 VDD.t465 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X89 VDD.t390 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 a_12612_160# VDD.t389 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X90 a_6034_296# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 term_2.t2 VSS.t536 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X91 vernier_delay_line_0.delay_unit_2_0.out_1.t5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X92 vernier_delay_line_0.start_neg.t1 diff_gen_0.delay_unit_2_6.in_1.t9 VSS.t158 VSS.t157 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X93 VSS.t40 start_buffer_0.start_buff.t12 diff_gen_0.delay_unit_2_1.in_2.t3 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X94 VDD.t148 diff_gen_0.delay_unit_2_5.in_2.t10 diff_gen_0.delay_unit_2_6.in_1.t5 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X95 VDD.t138 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X96 a_3364_2192.t1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 a_3628_2192.t3 VSS.t236 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X97 diff_gen_0.delay_unit_2_3.in_2.t5 diff_gen_0.delay_unit_2_2.in_1.t9 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X98 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X99 a_1346_2192.t5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 a_1082_2192.t1 VSS.t249 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X100 VDD.t283 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 VDD.t282 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X101 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 a_10474_2192.t5 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X102 VSS.t267 vernier_delay_line_0.stop_strong.t42 a_1082_2192.t6 VSS.t266 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X103 vernier_delay_line_0.stop_strong.t10 a_n6458_3464.t8 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X104 VDD.t51 diff_gen_0.delay_unit_2_4.in_1.t9 diff_gen_0.delay_unit_2_5.in_2.t0 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X105 a_14774_2192.t9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 a_14862_2192# VSS.t72 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X106 VSS.t544 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 VSS.t543 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X107 a_n6458_3464.t2 a_n6748_3464# VSS.t232 VSS.t231 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X108 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VDD.t221 VDD.t220 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X109 a_8732_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X110 VDD.t461 diff_gen_0.delay_unit_2_3.in_2.t9 diff_gen_0.delay_unit_2_3.in_1.t7 VDD.t460 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X111 VSS.t366 vernier_delay_line_0.stop_strong.t43 a_17056_2192.t11 VSS.t365 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X112 VDD.t435 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15162_730# VDD.t434 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X113 a_14774_2192.t0 vernier_delay_line_0.stop_strong.t44 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X114 a_5910_2192.t1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X115 a_n7038_3464# a_n7328_3464# VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X116 vernier_delay_line_0.delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 VSS.t318 VSS.t317 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X117 term_4.t0 a_10330_160# VSS.t483 VSS.t482 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X118 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VSS.t490 VSS.t489 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X119 a_10298_2192# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X120 VDD.t188 diff_gen_0.delay_unit_2_2.in_1.t10 diff_gen_0.delay_unit_2_2.in_2.t1 VDD.t187 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X121 VSS.t396 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 VSS.t395 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X122 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X123 VSS.t530 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 a_5766_160# VSS.t529 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X124 vernier_delay_line_0.stop_strong.t11 a_n6458_3464.t9 VSS.t123 VSS.t122 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X125 VDD.t453 vernier_delay_line_0.stop_strong.t45 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VDD.t452 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X126 a_4168_1376# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VSS.t344 VSS.t343 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X127 a_5646_2192.t3 vernier_delay_line_0.stop_strong.t46 VSS.t364 VSS.t363 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X128 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_11014_1376# a_10976_730# VDD.t491 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X129 a_17056_2192.t6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 a_17320_2192.t3 VSS.t75 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X130 VSS.t333 vernier_delay_line_0.stop_strong.t47 a_3364_2192.t4 VSS.t332 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X131 vernier_delay_line_0.stop_strong.t6 a_n6458_3464.t10 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X132 VSS.t287 diff_gen_0.delay_unit_2_4.in_2.t9 diff_gen_0.delay_unit_2_5.in_1.t2 VSS.t286 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X133 VSS.t467 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 VSS.t466 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X134 a_15038_2192.t3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 a_14774_2192.t3 VSS.t126 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X135 VDD.t430 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X136 a_6034_730# a_5766_160# term_2.t1 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X137 VDD.t293 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VDD.t292 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X138 a_n7038_3464# a_n7328_3464# VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X139 vernier_delay_line_0.start_pos.t3 diff_gen_0.delay_unit_2_6.in_2.t9 VSS.t192 VSS.t191 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X140 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X141 VSS.t510 a_13296_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VSS.t509 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X142 VSS.t128 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 VSS.t127 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X143 VSS.t257 vernier_delay_line_0.start_neg.t9 vernier_delay_line_0.start_pos.t0 VSS.t256 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X144 VSS.t448 diff_gen_0.delay_unit_2_3.in_1.t9 diff_gen_0.delay_unit_2_4.in_2.t2 VSS.t447 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X145 VDD.t144 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X146 VDD.t376 diff_gen_0.delay_unit_2_1.in_1.t9 diff_gen_0.delay_unit_2_1.in_2.t7 VDD.t375 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X147 VDD.t99 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X148 a_1346_2192.t1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X149 diff_gen_0.delay_unit_2_6.in_2.t6 diff_gen_0.delay_unit_2_5.in_1.t9 VDD.t335 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X150 VSS.t372 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 a_1202_160# VSS.t371 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X151 VSS.t316 diff_gen_0.delay_unit_2_2.in_2.t9 diff_gen_0.delay_unit_2_2.in_1.t6 VSS.t315 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X152 a_5734_2192# vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 a_5646_2192.t7 VSS.t463 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X153 diff_gen_0.delay_unit_2_6.in_2.t4 diff_gen_0.delay_unit_2_5.in_1.t10 VSS.t506 VSS.t505 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X154 a_8732_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X155 vernier_delay_line_0.stop_strong.t7 a_n6458_3464.t11 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X156 VDD.t186 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 VDD.t185 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X157 a_7928_2192.t8 vernier_delay_line_0.stop_strong.t48 VSS.t186 VSS.t185 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X158 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 vernier_delay_line_0.start_pos.t9 VDD.t480 VDD.t479 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X159 VSS.t277 vernier_delay_line_0.stop_strong.t49 a_5646_2192.t2 VSS.t276 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X160 VSS.t139 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 vernier_delay_line_0.delay_unit_2_0.out_1.t2 VSS.t138 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X161 VDD.t263 diff_gen_0.delay_unit_2_6.in_2.t10 diff_gen_0.delay_unit_2_6.in_1.t6 VDD.t262 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X162 vernier_delay_line_0.stop_strong.t8 a_n6458_3464.t12 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X163 VDD.t196 vernier_delay_line_0.stop_strong.t50 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X164 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 vernier_delay_line_0.stop_strong.t51 VDD.t250 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X165 diff_gen_0.delay_unit_2_3.in_1.t4 diff_gen_0.delay_unit_2_2.in_2.t10 VDD.t478 VDD.t477 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X166 term_4.t2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 VDD.t426 VDD.t425 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X167 vernier_delay_line_0.stop_strong.t9 a_n6458_3464.t13 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X168 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 a_5734_2192# VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X169 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VSS.t289 VSS.t288 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X170 VDD.t275 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 a_5766_160# VDD.t274 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X171 a_12492_2192.t1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 a_12756_2192.t3 VSS.t53 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X172 a_3452_2192# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X173 a_4168_1376# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VDD.t343 VDD.t342 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X174 a_n6748_3464# a_n7038_3464# VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X175 VSS.t213 vernier_delay_line_0.stop_strong.t52 a_10210_2192.t11 VSS.t212 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X176 diff_gen_0.delay_unit_2_2.in_2.t7 diff_gen_0.delay_unit_2_1.in_1.t10 VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X177 vernier_delay_line_0.delay_unit_2_0.out_1.t4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X178 a_12880_296# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 term_5.t2 VSS.t351 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X179 vernier_delay_line_0.stop_strong.t4 a_n6458_3464.t14 VSS.t96 VSS.t95 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X180 VDD.t497 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 VDD.t496 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X181 a_1170_2192# vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 a_1082_2192.t0 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X182 a_17860_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VSS.t379 VSS.t378 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X183 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 a_17320_2192.t5 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X184 VSS.t208 vernier_delay_line_0.stop_strong.t53 a_7928_2192.t7 VSS.t207 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X185 VDD.t396 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X186 diff_gen_0.delay_unit_2_2.in_1.t1 diff_gen_0.delay_unit_2_1.in_2.t10 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X187 VSS.t452 start_buffer_0.start_buff.t13 start_buffer_0.start_delay.t3 VSS.t451 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X188 VDD.t59 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X189 a_3364_2192.t9 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 a_3452_2192# VSS.t211 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X190 vernier_delay_line_0.stop_strong.t5 a_n6458_3464.t15 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X191 diff_gen_0.delay_unit_2_3.in_2.t4 diff_gen_0.delay_unit_2_2.in_1.t11 VDD.t457 VDD.t456 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X192 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 a_17822_296# VSS.t578 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X193 VDD.t71 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X194 VDD.t349 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 a_1202_160# VDD.t348 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X195 vernier_delay_line_0.stop_strong.t14 a_n6458_3464.t16 VSS.t200 VSS.t199 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X196 vernier_delay_line_0.stop_strong.t15 a_n6458_3464.t17 VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X197 a_12756_2192.t2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 a_12492_2192.t12 VSS.t174 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X198 VDD.t177 diff_gen_0.delay_unit_2_4.in_1.t10 diff_gen_0.delay_unit_2_4.in_2.t7 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X199 VDD.t404 diff_gen_0.delay_unit_2_6.in_1.t10 vernier_delay_line_0.start_neg.t5 VDD.t403 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X200 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 VSS.t146 VSS.t145 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X201 VDD.t493 vernier_delay_line_0.stop_strong.t54 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VDD.t492 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X202 VSS.t435 diff_gen_0.delay_unit_2_5.in_2.t11 diff_gen_0.delay_unit_2_5.in_1.t3 VSS.t434 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X203 a_n6748_3464# a_n7038_3464# VSS.t59 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X204 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 a_3628_2192.t5 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X205 term_1.t0 a_3484_160# VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X206 a_14774_2192.t2 vernier_delay_line_0.stop_strong.t55 VSS.t85 VSS.t84 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X207 a_17144_2192# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X208 vernier_delay_line_0.delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VSS.t320 VSS.t319 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X209 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 vernier_delay_line_0.stop_strong.t56 VDD.t232 VDD.t231 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X210 a_n7618_3464# a_n7908_3464# VDD.t241 VDD.t240 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X211 VSS.t398 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VSS.t397 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X212 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X213 VSS.t450 diff_gen_0.delay_unit_2_3.in_2.t10 diff_gen_0.delay_unit_2_4.in_1.t3 VSS.t449 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X214 a_5646_2192.t8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 a_5910_2192.t4 VSS.t566 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X215 vernier_delay_line_0.stop_strong.t30 a_n6458_3464.t18 VSS.t540 VSS.t539 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X216 VSS.t25 diff_gen_0.delay_unit_2_5.in_1.t11 diff_gen_0.delay_unit_2_6.in_2.t3 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X217 diff_gen_0.delay_unit_2_1.in_2.t2 start_buffer_0.start_buff.t14 VSS.t572 VSS.t571 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X218 a_8694_296# term_3.t4 VSS.t117 VSS.t116 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X219 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VDD.t449 VDD.t448 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X220 VSS.t465 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VSS.t464 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X221 VSS.t77 vernier_delay_line_0.stop_strong.t57 a_3364_2192.t3 VSS.t76 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X222 a_11014_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 VSS.t471 VSS.t470 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X223 vernier_delay_line_0.stop_strong.t31 a_n6458_3464.t19 VDD.t488 VDD.t487 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X224 vernier_delay_line_0.stop_strong.t2 a_n6458_3464.t20 VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X225 VDD.t39 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X226 a_1082_2192.t5 vernier_delay_line_0.stop_strong.t58 VSS.t293 VSS.t292 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X227 a_12880_730# a_12612_160# term_5.t1 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X228 a_17056_2192.t2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 a_17144_2192# VSS.t423 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X229 diff_gen_0.delay_unit_2_1.in_1.t4 start_buffer_0.start_delay.t10 VSS.t194 VSS.t193 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X230 VSS.t265 vernier_delay_line_0.start_pos.t10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VSS.t264 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X231 VSS.t368 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VSS.t367 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X232 a_17860_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X233 vernier_delay_line_0.stop_strong.t3 a_n6458_3464.t21 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X234 VDD.t217 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X235 VDD.t112 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X236 a_10210_2192.t2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 a_10474_2192.t3 VSS.t81 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X237 a_17056_2192.t10 vernier_delay_line_0.stop_strong.t59 VSS.t414 VSS.t413 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X238 a_8192_2192.t0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X239 VSS.t508 diff_gen_0.delay_unit_2_2.in_2.t11 diff_gen_0.delay_unit_2_3.in_1.t2 VSS.t507 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X240 VSS.t273 vernier_delay_line_0.start_neg.t10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 VSS.t272 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X241 a_n7618_3464# a_n7908_3464# VSS.t275 VSS.t274 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X242 diff_gen_0.delay_unit_2_5.in_1.t5 diff_gen_0.delay_unit_2_4.in_2.t10 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X243 VSS.t106 diff_gen_0.delay_unit_2_3.in_1.t10 diff_gen_0.delay_unit_2_3.in_2.t6 VSS.t105 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X244 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17860_1376# a_17822_730# VDD.t495 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X245 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X246 start_buffer_0.start_delay.t6 start_buffer_0.start_buff.t15 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X247 VSS.t210 a_1886_1376# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VSS.t209 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X248 VSS.t568 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 VSS.t567 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X249 a_n8488_3464# a_n8778_3464# VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X250 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 a_14862_2192# VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X251 a_5910_2192.t3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 a_5646_2192.t10 VSS.t255 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X252 VDD.t345 diff_gen_0.delay_unit_2_6.in_2.t11 vernier_delay_line_0.start_pos.t7 VDD.t344 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X253 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 vernier_delay_line_0.start_pos.t11 VDD.t211 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X254 a_8316_296# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 term_3.t0 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X255 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 VSS.t422 VSS.t421 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X256 VDD.t75 vernier_delay_line_0.stop_strong.t60 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X257 diff_gen_0.delay_unit_2_4.in_2.t5 diff_gen_0.delay_unit_2_3.in_1.t11 VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X258 a_7928_2192.t6 vernier_delay_line_0.stop_strong.t61 VSS.t552 VSS.t551 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X259 vernier_delay_line_0.stop_strong.t22 a_n6458_3464.t22 VSS.t327 VSS.t326 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X260 vernier_delay_line_0.stop_strong.t23 a_n6458_3464.t23 VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X261 term_1.t2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VDD.t226 VDD.t225 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X262 VSS.t497 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 VSS.t496 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X263 a_10298_2192# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 a_10210_2192.t7 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X264 vernier_delay_line_0.stop_strong.t28 a_n6458_3464.t24 VSS.t518 VSS.t517 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X265 VDD.t455 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X266 VSS.t165 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 a_8048_160# VSS.t164 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X267 term_7.t1 a_17176_160# VSS.t226 VSS.t225 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X268 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X269 a_8694_730# term_3.t5 VDD.t470 VDD.t469 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X270 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 a_1170_2192# VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X271 a_n6458_3464.t6 a_n6748_3464# VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X272 VSS.t52 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X273 start_buffer_0.start_delay.t2 start_buffer_0.start_buff.t16 VSS.t439 VSS.t438 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X274 a_11014_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VDD.t420 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X275 diff_gen_0.delay_unit_2_2.in_2.t6 diff_gen_0.delay_unit_2_1.in_1.t11 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X276 VSS.t431 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 VSS.t430 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X277 a_n8488_3464# a_n8778_3464# VSS.t446 VSS.t445 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X278 a_8016_2192# vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 a_7928_2192.t2 VSS.t524 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X279 start_buffer_0.start_buff.t7 a_n11872_5654# VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X280 VDD.t400 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VDD.t399 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X281 vernier_delay_line_0.stop_strong.t29 a_n6458_3464.t25 VSS.t520 VSS.t519 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X282 a_1346_2192.t4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 a_1082_2192.t3 VSS.t308 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X283 diff_gen_0.delay_unit_2_2.in_1.t2 diff_gen_0.delay_unit_2_1.in_2.t11 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X284 VSS.t101 diff_gen_0.delay_unit_2_4.in_2.t11 diff_gen_0.delay_unit_2_4.in_1.t0 VSS.t100 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X285 a_1848_296# term_0.t4 VSS.t196 VSS.t195 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X286 a_1470_296# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 term_0.t0 VSS.t493 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X287 vernier_delay_line_0.stop_strong.t24 a_n6458_3464.t26 VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X288 vernier_delay_line_0.delay_unit_2_0.out_1.t1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X289 VSS.t350 diff_gen_0.delay_unit_2_5.in_2.t12 diff_gen_0.delay_unit_2_6.in_1.t1 VSS.t349 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X290 VSS.t178 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10598_296# VSS.t177 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X291 VDD.t261 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VDD.t260 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X292 VSS.t481 vernier_delay_line_0.stop_strong.t62 a_12492_2192.t8 VSS.t480 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X293 diff_gen_0.delay_unit_2_3.in_2.t1 diff_gen_0.delay_unit_2_2.in_1.t12 VSS.t154 VSS.t153 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X294 diff_gen_0.delay_unit_2_1.in_2.t5 start_buffer_0.start_buff.t17 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X295 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 VSS.t83 VSS.t82 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X296 a_n6458_3464.t1 a_n6748_3464# VSS.t230 VSS.t229 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X297 VSS.t251 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VSS.t250 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X298 a_8316_730# a_8048_160# term_3.t3 VDD.t239 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X299 a_5734_2192# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X300 VSS.t548 diff_gen_0.delay_unit_2_4.in_1.t11 diff_gen_0.delay_unit_2_5.in_2.t6 VSS.t547 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X301 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 a_6412_296# VSS.t521 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X302 VSS.t171 vernier_delay_line_0.stop_strong.t63 a_12492_2192.t7 VSS.t170 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X303 VSS.t15 a_15578_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X304 a_5646_2192.t5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 a_5734_2192# VSS.t111 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X305 start_buffer_0.start_buff.t2 a_n11872_5654# VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X306 VSS.t137 diff_gen_0.delay_unit_2_3.in_2.t11 diff_gen_0.delay_unit_2_3.in_1.t6 VSS.t136 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X307 VDD.t386 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VDD.t385 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X308 a_3452_2192# vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 a_3364_2192.t8 VSS.t555 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X309 VDD.t142 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 a_8048_160# VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X310 term_7.t2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 VDD.t223 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X311 a_15540_296# term_6.t4 VSS.t119 VSS.t118 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X312 vernier_delay_line_0.stop_strong.t25 a_n6458_3464.t27 VSS.t362 VSS.t361 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X313 VDD.t394 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 vernier_delay_line_0.delay_unit_2_0.out_2 VDD.t393 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X314 diff_gen_0.delay_unit_2_4.in_1.t5 diff_gen_0.delay_unit_2_3.in_2.t12 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X315 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 VSS.t329 VSS.t328 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X316 a_17056_2192.t5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 a_17320_2192.t2 VSS.t47 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X317 VSS.t580 diff_gen_0.delay_unit_2_2.in_1.t13 diff_gen_0.delay_unit_2_2.in_2.t0 VSS.t579 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X318 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 VDD.t474 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X319 VSS.t224 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_6034_296# VSS.t223 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X320 a_1848_730# term_0.t5 VDD.t190 VDD.t189 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X321 a_1470_730# a_1202_160# term_0.t3 VDD.t251 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X322 diff_gen_0.delay_unit_2_5.in_1.t0 diff_gen_0.delay_unit_2_4.in_2.t12 VDD.t103 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X323 VSS.t374 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 VSS.t373 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X324 VDD.t155 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10598_730# VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X325 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X326 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VSS.t254 VSS.t253 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X327 a_3364_2192.t11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 a_3628_2192.t2 VSS.t299 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X328 VSS.t492 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 VSS.t491 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X329 VSS.t49 diff_gen_0.delay_unit_2_1.in_1.t12 diff_gen_0.delay_unit_2_1.in_2.t0 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X330 a_15162_296# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 term_6.t0 VSS.t386 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X331 diff_gen_0.delay_unit_2_6.in_2.t2 diff_gen_0.delay_unit_2_5.in_1.t12 VSS.t370 VSS.t369 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X332 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 vernier_delay_line_0.start_neg.t11 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X333 a_17144_2192# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 a_17056_2192.t1 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X334 diff_gen_0.delay_unit_2_4.in_2.t4 diff_gen_0.delay_unit_2_3.in_1.t12 VDD.t315 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X335 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_6450_1376# a_6412_730# VDD.t248 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X336 VSS.t306 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_3752_296# VSS.t305 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X337 VDD.t439 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VDD.t438 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X338 VSS.t526 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VSS.t525 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X339 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X340 a_10474_2192.t1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 a_10210_2192.t1 VSS.t415 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X341 VDD.t307 diff_gen_0.delay_unit_2_5.in_1.t13 diff_gen_0.delay_unit_2_5.in_2.t4 VDD.t306 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X342 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 vernier_delay_line_0.start_pos.t12 VSS.t218 VSS.t217 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X343 VDD.t327 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 VDD.t326 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X344 VSS.t535 diff_gen_0.delay_unit_2_6.in_2.t12 diff_gen_0.delay_unit_2_6.in_1.t7 VSS.t534 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X345 VSS.t244 a_8732_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VSS.t243 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X346 a_15540_730# term_6.t5 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X347 a_8192_2192.t3 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 a_7928_2192.t10 VSS.t575 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X348 diff_gen_0.delay_unit_2_3.in_1.t1 diff_gen_0.delay_unit_2_2.in_2.t12 VSS.t514 VSS.t513 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X349 diff_gen_0.delay_unit_2_1.in_1.t6 start_buffer_0.start_delay.t11 VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X350 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 vernier_delay_line_0.stop_strong.t64 VDD.t179 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X351 a_15038_2192.t1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X352 a_1170_2192# vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 a_1082_2192.t9 VSS.t356 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X353 a_8192_2192.t2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 a_7928_2192.t11 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X354 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X355 a_n11872_5654# start.t0 VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X356 diff_gen_0.delay_unit_2_2.in_2.t3 diff_gen_0.delay_unit_2_1.in_1.t13 VSS.t141 VSS.t140 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X357 VDD.t194 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_6034_730# VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X358 vernier_delay_line_0.delay_unit_2_0.out_1.t0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 VSS.t62 VSS.t61 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X359 VSS.t57 vernier_delay_line_0.stop_strong.t65 a_1082_2192.t4 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X360 VSS.t557 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VSS.t556 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X361 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VDD.t351 VDD.t350 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X362 VSS.t384 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 a_14894_160# VSS.t383 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X363 a_13296_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VSS.t113 VSS.t112 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X364 a_14774_2192.t8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 a_14862_2192# VSS.t252 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X365 diff_gen_0.delay_unit_2_2.in_1.t7 diff_gen_0.delay_unit_2_1.in_2.t12 VSS.t477 VSS.t476 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X366 diff_gen_0.delay_unit_2_3.in_2.t0 diff_gen_0.delay_unit_2_2.in_1.t14 VSS.t583 VSS.t582 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X367 VSS.t203 vernier_delay_line_0.stop_strong.t66 a_12492_2192.t6 VSS.t202 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X368 VSS.t454 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VSS.t453 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X369 a_15162_730# a_14894_160# term_6.t3 VDD.t368 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X370 VDD.t271 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_3752_730# VDD.t270 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X371 VDD.t57 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X372 VSS.t444 diff_gen_0.delay_unit_2_6.in_1.t11 vernier_delay_line_0.start_neg.t0 VSS.t443 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X373 diff_gen_0.delay_unit_2_6.in_1.t4 diff_gen_0.delay_unit_2_5.in_2.t13 VDD.t323 VDD.t322 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X374 VSS.t55 diff_gen_0.delay_unit_2_4.in_1.t12 diff_gen_0.delay_unit_2_4.in_2.t6 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X375 a_3628_2192.t1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 a_3364_2192.t0 VSS.t109 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X376 a_1082_2192.t10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 a_1170_2192# VSS.t296 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X377 VDD.t257 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 VDD.t256 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X378 VSS.t473 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 a_10330_160# VSS.t472 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X379 a_10474_2192.t4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X380 VDD.t311 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VDD.t310 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X381 a_n11872_5654# start.t1 VSS.t538 VSS.t537 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X382 VSS.t242 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17444_296# VSS.t241 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X383 VDD.t140 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDD.t139 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X384 diff_gen_0.delay_unit_2_5.in_2.t3 diff_gen_0.delay_unit_2_4.in_1.t13 VDD.t238 VDD.t237 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X385 a_14862_2192# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 a_14774_2192.t7 VSS.t455 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X386 VSS.t559 a_4168_1376# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VSS.t558 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X387 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 VSS.t64 VSS.t63 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X388 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 VDD.t464 VDD.t463 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X389 VSS.t504 vernier_delay_line_0.stop_strong.t67 a_14774_2192.t12 VSS.t503 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X390 vernier_delay_line_0.stop_strong.t26 a_n6458_3464.t28 VDD.t447 VDD.t446 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X391 VDD.t49 vernier_delay_line_0.stop_strong.t68 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X392 diff_gen_0.delay_unit_2_4.in_1.t4 diff_gen_0.delay_unit_2_3.in_2.t13 VDD.t353 VDD.t352 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X393 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VSS.t331 VSS.t330 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X394 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 vernier_delay_line_0.start_neg.t12 VDD.t269 VDD.t268 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X395 a_4130_296# term_1.t4 VSS.t259 VSS.t258 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X396 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 a_13258_296# VSS.t418 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X397 VDD.t367 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 a_14894_160# VDD.t366 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X398 a_12580_2192# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X399 VSS.t283 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 VSS.t282 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X400 a_13296_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VDD.t329 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X401 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X402 VDD.t41 start_buffer_0.start_delay.t12 diff_gen_0.delay_unit_2_1.in_1.t5 VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X403 VSS.t298 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 VSS.t297 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X404 a_5734_2192# vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 a_5646_2192.t12 VSS.t102 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X405 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X406 VSS.t546 vernier_delay_line_0.stop_strong.t69 a_5646_2192.t1 VSS.t545 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X407 a_3364_2192.t2 vernier_delay_line_0.stop_strong.t70 VSS.t74 VSS.t73 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X408 diff_gen_0.delay_unit_2_5.in_1.t7 diff_gen_0.delay_unit_2_4.in_2.t13 VSS.t533 VSS.t532 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X409 diff_gen_0.delay_unit_2_3.in_1.t3 diff_gen_0.delay_unit_2_2.in_2.t13 VDD.t273 VDD.t272 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X410 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 VSS.t459 VSS.t458 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X411 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 vernier_delay_line_0.stop_strong.t71 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X412 VSS.t169 vernier_delay_line_0.stop_strong.t72 a_17056_2192.t9 VSS.t168 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X413 a_12492_2192.t3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 a_12580_2192# VSS.t142 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X414 vernier_delay_line_0.stop_strong.t27 a_n6458_3464.t29 VSS.t502 VSS.t501 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X415 VSS.t475 diff_gen_0.delay_unit_2_6.in_2.t13 vernier_delay_line_0.start_pos.t2 VSS.t474 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X416 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 vernier_delay_line_0.start_pos.t13 VSS.t240 VSS.t239 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X417 VDD.t355 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 VDD.t354 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X418 diff_gen_0.delay_unit_2_4.in_2.t1 diff_gen_0.delay_unit_2_3.in_1.t13 VSS.t358 VSS.t357 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X419 VDD.t428 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 a_10330_160# VDD.t427 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X420 a_10298_2192# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 a_10210_2192.t6 VSS.t300 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X421 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VDD.t255 VDD.t254 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X422 VDD.t219 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17444_730# VDD.t218 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X423 a_3628_2192.t4 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X424 VDD.t398 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VDD.t397 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X425 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X426 term_5.t0 a_12612_160# VSS.t125 VSS.t124 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X427 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 a_12756_2192.t4 VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X428 VDD.t289 vernier_delay_line_0.start_pos.t14 vernier_delay_line_0.start_neg.t6 VDD.t288 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X429 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 VSS.t410 VSS.t409 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X430 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X431 a_6450_1376# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VSS.t420 VSS.t419 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X432 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X433 a_4130_730# term_1.t5 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X434 diff_gen_0.delay_unit_2_2.in_2.t2 diff_gen_0.delay_unit_2_1.in_1.t14 VSS.t94 VSS.t93 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X435 VDD.t357 diff_gen_0.delay_unit_2_6.in_1.t12 diff_gen_0.delay_unit_2_6.in_2.t1 VDD.t356 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X436 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13296_1376# a_13258_730# VDD.t462 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X437 a_17822_296# term_7.t4 VSS.t376 VSS.t375 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X438 VSS.t574 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 VSS.t573 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X439 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 VDD.t499 VDD.t498 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X440 a_12756_2192.t1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 a_12492_2192.t4 VSS.t201 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X441 a_n6458_3464.t5 a_n6748_3464# VDD.t201 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X442 diff_gen_0.delay_unit_2_2.in_1.t0 diff_gen_0.delay_unit_2_1.in_2.t13 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X443 VDD.t380 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 VDD.t379 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X444 a_10210_2192.t10 vernier_delay_line_0.stop_strong.t73 VSS.t360 VSS.t359 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X445 VDD.t484 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VDD.t483 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X446 VSS.t152 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 a_3484_160# VSS.t151 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X447 a_1886_1376# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VSS.t263 VSS.t262 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X448 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 vernier_delay_line_0.stop_strong.t74 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X449 diff_gen_0.delay_unit_2_6.in_1.t3 diff_gen_0.delay_unit_2_5.in_2.t14 VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X450 a_17320_2192.t4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X451 diff_gen_0.delay_unit_2_1.in_2.t1 start_buffer_0.start_buff.t18 VSS.t310 VSS.t309 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X452 a_3452_2192# vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 a_3364_2192.t7 VSS.t65 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X453 VDD.t114 diff_gen_0.delay_unit_2_2.in_1.t15 diff_gen_0.delay_unit_2_3.in_2.t3 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X454 a_1082_2192.t11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 a_1346_2192.t3 VSS.t498 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X455 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 VDD.t279 VDD.t278 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X456 vernier_delay_line_0.stop_strong.t0 a_n6458_3464.t30 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X457 VDD.t120 diff_gen_0.delay_unit_2_1.in_2.t14 diff_gen_0.delay_unit_2_1.in_1.t1 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X458 VDD.t95 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X459 vernier_delay_line_0.start_neg.t4 diff_gen_0.delay_unit_2_6.in_1.t13 VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X460 a_15038_2192.t2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 a_14774_2192.t4 VSS.t216 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X461 diff_gen_0.delay_unit_2_5.in_2.t1 diff_gen_0.delay_unit_2_4.in_1.t14 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X462 VSS.t295 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VSS.t294 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X463 VSS.t554 a_11014_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VSS.t553 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X464 VDD.t341 vernier_delay_line_0.stop_strong.t75 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VDD.t340 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X465 a_n6458_3464.t0 a_n6748_3464# VSS.t228 VSS.t227 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X466 term_5.t3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VDD.t392 VDD.t391 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X467 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 a_5910_2192.t0 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X468 VSS.t32 vernier_delay_line_0.stop_strong.t76 a_14774_2192.t1 VSS.t31 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X469 a_n7328_3464# a_n7618_3464# VDD.t163 VDD.t162 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X470 VSS.t130 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 vernier_delay_line_0.delay_unit_2_0.out_2 VSS.t129 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X471 a_6450_1376# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VDD.t445 VDD.t444 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X472 VDD.t77 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 VDD.t76 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X473 diff_gen_0.delay_unit_2_4.in_1.t2 diff_gen_0.delay_unit_2_3.in_2.t14 VSS.t402 VSS.t401 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X474 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X475 a_17822_730# term_7.t5 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X476 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 a_10298_2192# VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X477 VDD.t35 vernier_delay_line_0.stop_strong.t77 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X478 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 VSS.t512 VSS.t511 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X479 VDD.t173 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 VDD.t172 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X480 vernier_delay_line_0.stop_strong.t1 a_n6458_3464.t31 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X481 VSS.t34 vernier_delay_line_0.stop_strong.t78 a_5646_2192.t0 VSS.t33 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X482 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 vernier_delay_line_0.stop_strong.t79 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X483 term_3.t2 a_8048_160# VSS.t271 VSS.t270 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X484 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 a_8016_2192# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X485 a_17144_2192# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 a_17056_2192.t0 VSS.t131 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X486 diff_gen_0.delay_unit_2_5.in_1.t6 diff_gen_0.delay_unit_2_4.in_2.t14 VSS.t400 VSS.t399 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X487 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VSS.t461 VSS.t460 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X488 vernier_delay_line_0.stop_strong.t18 a_n6458_3464.t32 VDD.t265 VDD.t264 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X489 VDD.t136 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 a_3484_160# VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X490 a_1886_1376# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X491 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 VDD.t331 VDD.t330 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X492 a_10474_2192.t0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 a_10210_2192.t0 VSS.t78 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X493 VSS.t36 vernier_delay_line_0.stop_strong.t80 a_17056_2192.t8 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X494 a_10976_296# term_4.t4 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X495 a_n7328_3464# a_n7618_3464# VSS.t184 VSS.t183 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X496 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 vernier_delay_line_0.start_neg.t13 VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X497 start_buffer_0.start_delay.t5 start_buffer_0.start_buff.t19 VDD.t277 VDD.t276 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X498 diff_gen_0.delay_unit_2_4.in_2.t0 diff_gen_0.delay_unit_2_3.in_1.t14 VSS.t285 VSS.t284 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X499 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X500 VSS.t442 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 a_17176_160# VSS.t441 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X501 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 a_1346_2192.t0 VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X502 term_2.t0 a_5766_160# VSS.t173 VSS.t172 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X503 a_n8198_3464# a_n8488_3464# VDD.t285 VDD.t284 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X504 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VSS.t408 VSS.t407 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X505 vernier_delay_line_0.start_pos.t6 diff_gen_0.delay_unit_2_6.in_2.t14 VDD.t418 VDD.t417 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X506 VSS.t215 diff_gen_0.delay_unit_2_5.in_1.t14 diff_gen_0.delay_unit_2_5.in_2.t2 VSS.t214 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X507 VDD.t422 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VDD.t421 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X508 a_14862_2192# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 VSS.t382 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X509 a_5646_2192.t6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 a_5734_2192# VSS.t462 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X510 VSS.t71 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VSS.t70 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X511 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X512 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X513 vernier_delay_line_0.stop_strong.t19 a_n6458_3464.t33 VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X514 VSS.t38 vernier_delay_line_0.stop_strong.t81 a_7928_2192.t5 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X515 diff_gen_0.delay_unit_2_1.in_1.t3 start_buffer_0.start_delay.t13 VSS.t323 VSS.t322 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X516 a_12580_2192# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 a_12492_2192.t10 VSS.t235 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X517 vernier_delay_line_0.stop_strong.t20 a_n6458_3464.t34 VSS.t325 VSS.t324 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X518 VDD.t230 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VDD.t229 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X519 a_10210_2192.t9 vernier_delay_line_0.stop_strong.t82 VSS.t302 VSS.t301 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X520 vernier_delay_line_0.stop_strong.t21 a_n6458_3464.t35 VDD.t303 VDD.t302 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X521 term_0.t2 a_1202_160# VSS.t281 VSS.t280 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X522 a_10598_296# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 term_4.t3 VSS.t469 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X523 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 a_3452_2192# VSS.t86 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X524 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 VSS.t404 VSS.t403 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X525 start_buffer_0.start_delay.t1 start_buffer_0.start_buff.t20 VSS.t433 VSS.t432 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X526 a_12580_2192# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 a_12492_2192.t2 VSS.t97 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X527 term_3.t1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X528 a_n8198_3464# a_n8488_3464# VSS.t314 VSS.t313 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X529 VDD.t374 diff_gen_0.delay_unit_2_1.in_1.t15 diff_gen_0.delay_unit_2_2.in_2.t5 VDD.t373 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X530 start_buffer_0.start_buff.t6 a_n11872_5654# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X531 a_6412_296# term_2.t4 VSS.t495 VSS.t494 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X532 VDD.t468 start_buffer_0.start_delay.t14 start_buffer_0.start_buff.t9 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X533 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X534 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 a_15540_296# VSS.t381 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X535 vernier_delay_line_0.stop_strong.t12 a_n6458_3464.t36 VSS.t198 VSS.t197 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X536 VDD.t209 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VDD.t208 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X537 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 a_15038_2192.t0 VSS.t385 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X538 VDD.t171 diff_gen_0.delay_unit_2_1.in_2.t15 diff_gen_0.delay_unit_2_2.in_1.t3 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X539 a_10976_730# term_4.t5 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X540 a_3628_2192.t0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 a_3364_2192.t12 VSS.t110 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X541 vernier_delay_line_0.stop_strong.t13 a_n6458_3464.t37 VDD.t167 VDD.t166 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X542 VSS.t205 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 VSS.t204 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X543 diff_gen_0.delay_unit_2_6.in_1.t0 diff_gen_0.delay_unit_2_5.in_2.t15 VSS.t115 VSS.t114 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X544 VDD.t406 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 a_17176_160# VDD.t405 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X545 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X546 term_2.t3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VDD.t459 VDD.t458 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X547 a_12492_2192.t11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 a_12756_2192.t0 VSS.t321 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X548 a_8016_2192# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VSS.t162 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X549 vernier_delay_line_0.stop_strong.t16 a_n6458_3464.t38 VSS.t220 VSS.t219 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X550 VDD.t441 start_buffer_0.start_buff.t21 diff_gen_0.delay_unit_2_1.in_2.t4 VDD.t440 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X551 vernier_delay_line_0.start_neg.t3 diff_gen_0.delay_unit_2_6.in_1.t14 VDD.t321 VDD.t320 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X552 VSS.t80 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 VSS.t79 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X553 VSS.t304 vernier_delay_line_0.stop_strong.t83 a_14774_2192.t5 VSS.t303 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X554 VSS.t340 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 VSS.t339 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X555 diff_gen_0.delay_unit_2_5.in_2.t5 diff_gen_0.delay_unit_2_4.in_1.t15 VSS.t406 VSS.t405 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X556 a_12492_2192.t5 vernier_delay_line_0.stop_strong.t84 VSS.t238 VSS.t237 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X557 start_buffer_0.start_buff.t1 a_n11872_5654# VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X558 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 a_17144_2192# VSS.t440 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X559 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 VSS.t394 VSS.t393 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X560 VDD.t378 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VDD.t377 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X561 a_n7908_3464# a_n8198_3464# VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X562 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 vernier_delay_line_0.stop_strong.t85 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X563 diff_gen_0.delay_unit_2_4.in_1.t1 diff_gen_0.delay_unit_2_3.in_2.t15 VSS.t528 VSS.t527 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X564 term_0.t1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X565 a_10598_730# a_10330_160# term_4.t1 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X566 a_17320_2192.t1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 a_17056_2192.t7 VSS.t206 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X567 vernier_delay_line_0.stop_strong.t17 a_n6458_3464.t39 VSS.t222 VSS.t221 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X568 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 vernier_delay_line_0.start_neg.t14 VSS.t479 VSS.t478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X569 vernier_delay_line_0.delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X570 start_buffer_0.start_delay.t4 start_buffer_0.start_buff.t22 VDD.t476 VDD.t475 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X571 term_6.t2 a_14894_160# VSS.t390 VSS.t389 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X572 a_17320_2192.t0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 a_17056_2192.t4 VSS.t377 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X573 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X574 VSS.t500 start_buffer_0.start_delay.t15 diff_gen_0.delay_unit_2_1.in_1.t2 VSS.t499 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X575 a_6412_730# term_2.t5 VDD.t287 VDD.t286 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X576 a_3752_296# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 term_1.t3 VSS.t107 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X577 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 VSS.t269 VSS.t268 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X578 VSS.t412 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12880_296# VSS.t411 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X579 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15578_1376# a_15540_730# VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X580 VDD.t372 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 VDD.t371 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X581 VSS.t246 vernier_delay_line_0.stop_strong.t86 a_10210_2192.t8 VSS.t245 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X582 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 a_8192_2192.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X583 diff_gen_0.delay_unit_2_3.in_1.t0 diff_gen_0.delay_unit_2_2.in_2.t14 VSS.t429 VSS.t428 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X584 VDD.t243 diff_gen_0.delay_unit_2_4.in_2.t15 diff_gen_0.delay_unit_2_5.in_1.t1 VDD.t242 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X585 a_n7908_3464# a_n8198_3464# VSS.t144 VSS.t143 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X586 VDD.t412 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 VDD.t411 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X587 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 a_8694_296# VSS.t161 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X588 VSS.t565 a_17860_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VSS.t564 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X589 VSS.t248 vernier_delay_line_0.stop_strong.t87 a_7928_2192.t4 VSS.t247 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X590 start_buffer_0.start_buff.t5 a_n11872_5654# VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X591 VSS.t182 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 VSS.t181 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X592 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 a_12580_2192# VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X593 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 VSS.t487 VSS.t486 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X594 a_5646_2192.t11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 a_5910_2192.t2 VSS.t26 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X595 a_n8778_3464# stop.t0 VDD.t161 VDD.t160 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X596 vernier_delay_line_0.start_pos.t5 diff_gen_0.delay_unit_2_6.in_2.t15 VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X597 VDD.t65 vernier_delay_line_0.start_neg.t15 vernier_delay_line_0.start_pos.t1 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X598 VDD.t236 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 VDD.t235 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X599 VDD.t67 diff_gen_0.delay_unit_2_3.in_1.t15 diff_gen_0.delay_unit_2_4.in_2.t3 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X600 start_buffer_0.start_delay.t0 start_buffer_0.start_buff.t23 VSS.t425 VSS.t424 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X601 VDD.t245 diff_gen_0.delay_unit_2_2.in_2.t15 diff_gen_0.delay_unit_2_2.in_1.t4 VDD.t244 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X602 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VSS.t160 VSS.t159 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X603 a_10210_2192.t5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 a_10298_2192# VSS.t108 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X604 diff_gen_0.delay_unit_2_6.in_2.t5 diff_gen_0.delay_unit_2_5.in_1.t15 VDD.t207 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X605 VSS.t561 vernier_delay_line_0.start_pos.t15 vernier_delay_line_0.start_neg.t7 VSS.t560 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X606 a_10210_2192.t4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 a_10298_2192# VSS.t522 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X607 a_7928_2192.t1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 a_8016_2192# VSS.t163 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X608 VDD.t490 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 vernier_delay_line_0.delay_unit_2_0.out_1.t3 VDD.t489 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X609 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 VSS.t99 VSS.t98 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X610 a_n6458_3464.t4 a_n6748_3464# VDD.t199 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X611 VSS.t167 diff_gen_0.delay_unit_2_6.in_1.t15 diff_gen_0.delay_unit_2_6.in_2.t0 VSS.t166 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X612 VSS.t417 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8316_296# VSS.t416 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X613 start_buffer_0.start_buff.t0 a_n11872_5654# VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X614 term_6.t1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VDD.t361 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X615 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VSS.t577 VSS.t576 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.15
X616 a_3752_730# a_3484_160# term_1.t1 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X617 a_7928_2192.t0 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 a_8016_2192# VSS.t523 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X618 a_n8778_3464# stop.t1 VSS.t516 VSS.t515 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X619 VSS.t392 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VSS.t391 sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X620 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 VDD.t501 VDD.t500 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X621 VDD.t384 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12880_730# VDD.t383 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X622 start_buffer_0.start_buff.t4 a_n11872_5654# VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
X623 a_1082_2192.t2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 a_1346_2192.t2 VSS.t307 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
R0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 890.727
R1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 742.783
R2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 665.16
R3 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 623.388
R4 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 523.774
R5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 431.807
R6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 427.875
R7 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 364.733
R8 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 208.5
R9 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 168.007
R10 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 75.2663
R11 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 31.2728
R12 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 31.0337
R13 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 9.52217
R14 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R15 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 9.08234
R16 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R17 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 4.50239
R18 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 0.898227
R19 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 0.707022
R20 VDD.n926 VDD.n72 2106.47
R21 VDD.n940 VDD.n64 2106.47
R22 VDD.n954 VDD.n56 2106.47
R23 VDD.n968 VDD.n48 2106.47
R24 VDD.n982 VDD.n40 2106.47
R25 VDD.n996 VDD.n32 2106.47
R26 VDD.n1010 VDD.n24 2106.47
R27 VDD.n13 VDD.n7 2106.47
R28 VDD.n930 VDD.n925 2101.76
R29 VDD.n944 VDD.n939 2101.76
R30 VDD.n958 VDD.n953 2101.76
R31 VDD.n972 VDD.n967 2101.76
R32 VDD.n986 VDD.n981 2101.76
R33 VDD.n1000 VDD.n995 2101.76
R34 VDD.n1014 VDD.n1009 2101.76
R35 VDD.n9 VDD.n8 2101.76
R36 VDD.n910 VDD.n721 2093.75
R37 VDD.n895 VDD.n729 2093.75
R38 VDD.n880 VDD.n737 2093.75
R39 VDD.n865 VDD.n745 2093.75
R40 VDD.n850 VDD.n753 2093.75
R41 VDD.n835 VDD.n761 2093.75
R42 VDD.n820 VDD.n769 2093.75
R43 VDD.n805 VDD.n777 2093.75
R44 VDD.n790 VDD.n785 2093.75
R45 VDD.n650 VDD.n548 2093.75
R46 VDD.n661 VDD.n535 2093.75
R47 VDD.n672 VDD.n522 2093.75
R48 VDD.n683 VDD.n509 2093.75
R49 VDD.n694 VDD.n496 2093.75
R50 VDD.n705 VDD.n483 2093.75
R51 VDD.n479 VDD.n478 2093.75
R52 VDD.n915 VDD.n722 2088.75
R53 VDD.n900 VDD.n730 2088.75
R54 VDD.n885 VDD.n738 2088.75
R55 VDD.n870 VDD.n746 2088.75
R56 VDD.n855 VDD.n754 2088.75
R57 VDD.n840 VDD.n762 2088.75
R58 VDD.n825 VDD.n770 2088.75
R59 VDD.n810 VDD.n778 2088.75
R60 VDD.n795 VDD.n786 2088.75
R61 VDD.n642 VDD.n554 2088.75
R62 VDD.n653 VDD.n541 2088.75
R63 VDD.n664 VDD.n528 2088.75
R64 VDD.n675 VDD.n515 2088.75
R65 VDD.n686 VDD.n502 2088.75
R66 VDD.n697 VDD.n489 2088.75
R67 VDD.n708 VDD.n474 2088.75
R68 VDD.n461 VDD.n459 1643.42
R69 VDD.n451 VDD.n449 1643.42
R70 VDD.n441 VDD.n439 1643.42
R71 VDD.n431 VDD.n429 1643.42
R72 VDD.n421 VDD.n419 1643.42
R73 VDD.n411 VDD.n409 1643.42
R74 VDD.n401 VDD.n399 1643.42
R75 VDD.n392 VDD.n390 1643.42
R76 VDD.n459 VDD.n458 1586.75
R77 VDD.n449 VDD.n448 1586.75
R78 VDD.n439 VDD.n438 1586.75
R79 VDD.n429 VDD.n428 1586.75
R80 VDD.n419 VDD.n418 1586.75
R81 VDD.n409 VDD.n408 1586.75
R82 VDD.n399 VDD.n398 1586.75
R83 VDD.n390 VDD.n389 1586.75
R84 VDD.n928 VDD.n925 1450
R85 VDD.n942 VDD.n939 1450
R86 VDD.n956 VDD.n953 1450
R87 VDD.n970 VDD.n967 1450
R88 VDD.n984 VDD.n981 1450
R89 VDD.n998 VDD.n995 1450
R90 VDD.n1012 VDD.n1009 1450
R91 VDD.n10 VDD.n8 1450
R92 VDD.n911 VDD.n721 1326.32
R93 VDD.n896 VDD.n729 1326.32
R94 VDD.n881 VDD.n737 1326.32
R95 VDD.n866 VDD.n745 1326.32
R96 VDD.n851 VDD.n753 1326.32
R97 VDD.n836 VDD.n761 1326.32
R98 VDD.n821 VDD.n769 1326.32
R99 VDD.n806 VDD.n777 1326.32
R100 VDD.n791 VDD.n785 1326.32
R101 VDD.n638 VDD.n548 1326.32
R102 VDD.n545 VDD.n535 1326.32
R103 VDD.n532 VDD.n522 1326.32
R104 VDD.n519 VDD.n509 1326.32
R105 VDD.n506 VDD.n496 1326.32
R106 VDD.n493 VDD.n483 1326.32
R107 VDD.n480 VDD.n479 1326.32
R108 VDD.n181 VDD.n180 1126.67
R109 VDD.n184 VDD.n183 1126.67
R110 VDD.n187 VDD.n186 1126.67
R111 VDD.n190 VDD.n189 1126.67
R112 VDD.n193 VDD.n192 1126.67
R113 VDD.n196 VDD.n195 1126.67
R114 VDD.n199 VDD.n198 1126.67
R115 VDD.n202 VDD.n201 1126.67
R116 VDD.n205 VDD.n204 1126.67
R117 VDD.n208 VDD.n207 1126.67
R118 VDD.n211 VDD.n210 1126.67
R119 VDD.n214 VDD.n213 1126.67
R120 VDD.n217 VDD.n216 1126.67
R121 VDD.n220 VDD.n219 1126.67
R122 VDD.n223 VDD.n222 1126.67
R123 VDD.n226 VDD.n225 1126.67
R124 VDD.n229 VDD.n228 1126.67
R125 VDD.n232 VDD.n231 1126.67
R126 VDD.n235 VDD.n234 1126.67
R127 VDD.n238 VDD.n237 1126.67
R128 VDD.n241 VDD.n240 1126.67
R129 VDD.n244 VDD.n243 1126.67
R130 VDD.n247 VDD.n246 1126.67
R131 VDD.n250 VDD.n249 1126.67
R132 VDD.n253 VDD.n252 1126.67
R133 VDD.n178 VDD.n177 1126.67
R134 VDD.n175 VDD.n174 1126.67
R135 VDD.n591 VDD.n590 1126.67
R136 VDD.n594 VDD.n593 1126.67
R137 VDD.n597 VDD.n596 1126.67
R138 VDD.n600 VDD.n599 1126.67
R139 VDD.n603 VDD.n602 1126.67
R140 VDD.n588 VDD.n587 1126.67
R141 VDD.n585 VDD.n584 1126.67
R142 VDD.n933 VDD.n69 224.69
R143 VDD.n947 VDD.n61 224.69
R144 VDD.n961 VDD.n53 224.69
R145 VDD.n975 VDD.n45 224.69
R146 VDD.n989 VDD.n37 224.69
R147 VDD.n1003 VDD.n29 224.69
R148 VDD.n1017 VDD.n21 224.69
R149 VDD.n15 VDD.n6 224.69
R150 VDD.n932 VDD.n931 224.189
R151 VDD.n946 VDD.n945 224.189
R152 VDD.n960 VDD.n959 224.189
R153 VDD.n974 VDD.n973 224.189
R154 VDD.n988 VDD.n987 224.189
R155 VDD.n1002 VDD.n1001 224.189
R156 VDD.n1016 VDD.n1015 224.189
R157 VDD.n14 VDD.n0 224.189
R158 VDD.n909 VDD.n720 223.333
R159 VDD.n894 VDD.n728 223.333
R160 VDD.n879 VDD.n736 223.333
R161 VDD.n864 VDD.n744 223.333
R162 VDD.n849 VDD.n752 223.333
R163 VDD.n834 VDD.n760 223.333
R164 VDD.n819 VDD.n768 223.333
R165 VDD.n804 VDD.n776 223.333
R166 VDD.n789 VDD.n784 223.333
R167 VDD.n649 VDD.n549 223.333
R168 VDD.n660 VDD.n536 223.333
R169 VDD.n671 VDD.n523 223.333
R170 VDD.n682 VDD.n510 223.333
R171 VDD.n693 VDD.n497 223.333
R172 VDD.n704 VDD.n484 223.333
R173 VDD.n473 VDD.n468 223.333
R174 VDD.n916 VDD.n715 222.8
R175 VDD.n901 VDD.n723 222.8
R176 VDD.n886 VDD.n731 222.8
R177 VDD.n871 VDD.n739 222.8
R178 VDD.n856 VDD.n747 222.8
R179 VDD.n841 VDD.n755 222.8
R180 VDD.n826 VDD.n763 222.8
R181 VDD.n811 VDD.n771 222.8
R182 VDD.n796 VDD.n779 222.8
R183 VDD.n644 VDD.n643 222.8
R184 VDD.n655 VDD.n654 222.8
R185 VDD.n666 VDD.n665 222.8
R186 VDD.n677 VDD.n676 222.8
R187 VDD.n688 VDD.n687 222.8
R188 VDD.n699 VDD.n698 222.8
R189 VDD.n710 VDD.n709 222.8
R190 VDD.n462 VDD.t208 196.429
R191 VDD.n452 VDD.t395 196.429
R192 VDD.n442 VDD.t483 196.429
R193 VDD.n432 VDD.t143 196.429
R194 VDD.n422 VDD.t429 196.429
R195 VDD.n412 VDD.t454 196.429
R196 VDD.n402 VDD.t229 196.429
R197 VDD.n393 VDD.t38 196.429
R198 VDD.n464 VDD.n458 184.671
R199 VDD.n454 VDD.n448 184.671
R200 VDD.n444 VDD.n438 184.671
R201 VDD.n434 VDD.n428 184.671
R202 VDD.n424 VDD.n418 184.671
R203 VDD.n414 VDD.n408 184.671
R204 VDD.n404 VDD.n398 184.671
R205 VDD.n395 VDD.n389 184.671
R206 VDD.n460 VDD.t131 183.929
R207 VDD.n450 VDD.t150 183.929
R208 VDD.n440 VDD.t227 183.929
R209 VDD.n430 VDD.t2 183.929
R210 VDD.n420 VDD.t415 183.929
R211 VDD.n410 VDD.t350 183.929
R212 VDD.n400 VDD.t364 183.929
R213 VDD.n391 VDD.t220 183.929
R214 VDD.n174 VDD.n79 181.25
R215 VDD.n174 VDD.n81 181.25
R216 VDD.n177 VDD.n81 181.25
R217 VDD.n177 VDD.n86 181.25
R218 VDD.n180 VDD.n86 181.25
R219 VDD.n180 VDD.n88 181.25
R220 VDD.n183 VDD.n88 181.25
R221 VDD.n183 VDD.n93 181.25
R222 VDD.n186 VDD.n93 181.25
R223 VDD.n186 VDD.n95 181.25
R224 VDD.n189 VDD.n95 181.25
R225 VDD.n189 VDD.n100 181.25
R226 VDD.n192 VDD.n100 181.25
R227 VDD.n192 VDD.n102 181.25
R228 VDD.n195 VDD.n102 181.25
R229 VDD.n195 VDD.n107 181.25
R230 VDD.n198 VDD.n107 181.25
R231 VDD.n198 VDD.n109 181.25
R232 VDD.n201 VDD.n109 181.25
R233 VDD.n201 VDD.n114 181.25
R234 VDD.n204 VDD.n114 181.25
R235 VDD.n204 VDD.n116 181.25
R236 VDD.n207 VDD.n116 181.25
R237 VDD.n207 VDD.n121 181.25
R238 VDD.n210 VDD.n121 181.25
R239 VDD.n210 VDD.n123 181.25
R240 VDD.n213 VDD.n123 181.25
R241 VDD.n213 VDD.n128 181.25
R242 VDD.n216 VDD.n128 181.25
R243 VDD.n216 VDD.n130 181.25
R244 VDD.n219 VDD.n130 181.25
R245 VDD.n219 VDD.n135 181.25
R246 VDD.n222 VDD.n135 181.25
R247 VDD.n222 VDD.n137 181.25
R248 VDD.n225 VDD.n137 181.25
R249 VDD.n225 VDD.n142 181.25
R250 VDD.n228 VDD.n142 181.25
R251 VDD.n228 VDD.n144 181.25
R252 VDD.n231 VDD.n144 181.25
R253 VDD.n231 VDD.n149 181.25
R254 VDD.n234 VDD.n149 181.25
R255 VDD.n234 VDD.n151 181.25
R256 VDD.n237 VDD.n151 181.25
R257 VDD.n237 VDD.n156 181.25
R258 VDD.n240 VDD.n156 181.25
R259 VDD.n240 VDD.n158 181.25
R260 VDD.n243 VDD.n158 181.25
R261 VDD.n243 VDD.n163 181.25
R262 VDD.n246 VDD.n163 181.25
R263 VDD.n246 VDD.n165 181.25
R264 VDD.n249 VDD.n165 181.25
R265 VDD.n249 VDD.n170 181.25
R266 VDD.n252 VDD.n170 181.25
R267 VDD.n252 VDD.n172 181.25
R268 VDD.n584 VDD.n559 181.25
R269 VDD.n584 VDD.n561 181.25
R270 VDD.n587 VDD.n561 181.25
R271 VDD.n587 VDD.n566 181.25
R272 VDD.n590 VDD.n566 181.25
R273 VDD.n590 VDD.n568 181.25
R274 VDD.n593 VDD.n568 181.25
R275 VDD.n593 VDD.n573 181.25
R276 VDD.n596 VDD.n573 181.25
R277 VDD.n596 VDD.n575 181.25
R278 VDD.n599 VDD.n575 181.25
R279 VDD.n599 VDD.n580 181.25
R280 VDD.n602 VDD.n580 181.25
R281 VDD.n602 VDD.n582 181.25
R282 VDD.n464 VDD.n357 175.298
R283 VDD.n454 VDD.n361 175.298
R284 VDD.n444 VDD.n365 175.298
R285 VDD.n434 VDD.n369 175.298
R286 VDD.n424 VDD.n373 175.298
R287 VDD.n414 VDD.n377 175.298
R288 VDD.n404 VDD.n381 175.298
R289 VDD.n395 VDD.n385 175.298
R290 VDD.n256 VDD.n255 175.123
R291 VDD.n173 VDD.n77 175.123
R292 VDD.n606 VDD.n605 175.123
R293 VDD.n583 VDD.n557 175.123
R294 VDD.t296 VDD.n926 169.983
R295 VDD.t342 VDD.n940 169.983
R296 VDD.t444 VDD.n954 169.983
R297 VDD.t0 VDD.n968 169.983
R298 VDD.t419 VDD.n982 169.983
R299 VDD.t328 VDD.n996 169.983
R300 VDD.t362 VDD.n1010 169.983
R301 VDD.t86 VDD.n7 169.983
R302 VDD.n930 VDD.t348 164.046
R303 VDD.n944 VDD.t135 164.046
R304 VDD.n958 VDD.t274 164.046
R305 VDD.n972 VDD.t141 164.046
R306 VDD.n986 VDD.t427 164.046
R307 VDD.n1000 VDD.t389 164.046
R308 VDD.n1014 VDD.t366 164.046
R309 VDD.t405 VDD.n9 164.046
R310 VDD.n176 VDD.t446 160.923
R311 VDD.t90 VDD.n176 160.923
R312 VDD.n179 VDD.t90 160.923
R313 VDD.t266 VDD.n179 160.923
R314 VDD.n182 VDD.t266 160.923
R315 VDD.t304 VDD.n182 160.923
R316 VDD.n185 VDD.t304 160.923
R317 VDD.t84 VDD.n185 160.923
R318 VDD.n188 VDD.t84 160.923
R319 VDD.t166 VDD.n188 160.923
R320 VDD.n191 VDD.t166 160.923
R321 VDD.t332 VDD.n191 160.923
R322 VDD.n194 VDD.t332 160.923
R323 VDD.t487 VDD.n194 160.923
R324 VDD.n197 VDD.t487 160.923
R325 VDD.t108 VDD.n197 160.923
R326 VDD.n200 VDD.t108 160.923
R327 VDD.t6 VDD.n200 160.923
R328 VDD.n203 VDD.t6 160.923
R329 VDD.t168 VDD.n203 160.923
R330 VDD.n206 VDD.t168 160.923
R331 VDD.t88 VDD.n206 160.923
R332 VDD.n209 VDD.t88 160.923
R333 VDD.t264 VDD.n209 160.923
R334 VDD.n212 VDD.t264 160.923
R335 VDD.t42 VDD.n212 160.923
R336 VDD.n215 VDD.t42 160.923
R337 VDD.t106 VDD.n215 160.923
R338 VDD.n218 VDD.t106 160.923
R339 VDD.t302 VDD.n218 160.923
R340 VDD.n221 VDD.t302 160.923
R341 VDD.t202 VDD.n221 160.923
R342 VDD.n224 VDD.t202 160.923
R343 VDD.t198 VDD.n224 160.923
R344 VDD.n227 VDD.t198 160.923
R345 VDD.t204 VDD.n227 160.923
R346 VDD.n230 VDD.t204 160.923
R347 VDD.t200 VDD.n230 160.923
R348 VDD.n233 VDD.t200 160.923
R349 VDD.t52 VDD.n233 160.923
R350 VDD.n236 VDD.t52 160.923
R351 VDD.t13 VDD.n236 160.923
R352 VDD.n239 VDD.t13 160.923
R353 VDD.t162 VDD.n239 160.923
R354 VDD.n242 VDD.t162 160.923
R355 VDD.t240 VDD.n242 160.923
R356 VDD.n245 VDD.t240 160.923
R357 VDD.t123 VDD.n245 160.923
R358 VDD.n248 VDD.t123 160.923
R359 VDD.t284 VDD.n248 160.923
R360 VDD.n251 VDD.t284 160.923
R361 VDD.t407 VDD.n251 160.923
R362 VDD.n254 VDD.t407 160.923
R363 VDD.t160 VDD.n254 160.923
R364 VDD.n586 VDD.t475 160.923
R365 VDD.t276 VDD.n586 160.923
R366 VDD.n589 VDD.t276 160.923
R367 VDD.t68 VDD.n589 160.923
R368 VDD.n592 VDD.t68 160.923
R369 VDD.t18 VDD.n592 160.923
R370 VDD.n595 VDD.t18 160.923
R371 VDD.t20 VDD.n595 160.923
R372 VDD.n598 VDD.t20 160.923
R373 VDD.t22 VDD.n598 160.923
R374 VDD.n601 VDD.t22 160.923
R375 VDD.t16 VDD.n601 160.923
R376 VDD.n604 VDD.t16 160.923
R377 VDD.t191 VDD.n604 160.923
R378 VDD.n911 VDD.n720 158.292
R379 VDD.n896 VDD.n728 158.292
R380 VDD.n881 VDD.n736 158.292
R381 VDD.n866 VDD.n744 158.292
R382 VDD.n851 VDD.n752 158.292
R383 VDD.n836 VDD.n760 158.292
R384 VDD.n821 VDD.n768 158.292
R385 VDD.n806 VDD.n776 158.292
R386 VDD.n791 VDD.n784 158.292
R387 VDD.n638 VDD.n549 158.292
R388 VDD.n545 VDD.n536 158.292
R389 VDD.n532 VDD.n523 158.292
R390 VDD.n519 VDD.n510 158.292
R391 VDD.n506 VDD.n497 158.292
R392 VDD.n493 VDD.n484 158.292
R393 VDD.n480 VDD.n473 158.292
R394 VDD.n932 VDD.n73 154.667
R395 VDD.n946 VDD.n65 154.667
R396 VDD.n960 VDD.n57 154.667
R397 VDD.n974 VDD.n49 154.667
R398 VDD.n988 VDD.n41 154.667
R399 VDD.n1002 VDD.n33 154.667
R400 VDD.n1016 VDD.n25 154.667
R401 VDD.n14 VDD.n2 154.667
R402 VDD.t210 VDD.n910 151.868
R403 VDD.t369 VDD.n895 151.868
R404 VDD.t181 VDD.n880 151.868
R405 VDD.t481 VDD.n865 151.868
R406 VDD.t473 VDD.n850 151.868
R407 VDD.t298 VDD.n835 151.868
R408 VDD.t92 VDD.n820 151.868
R409 VDD.t280 VDD.n805 151.868
R410 VDD.t409 VDD.n790 151.868
R411 VDD.n478 VDD.t145 151.868
R412 VDD.t178 VDD.n461 146.282
R413 VDD.t26 VDD.n451 146.282
R414 VDD.t214 VDD.n441 146.282
R415 VDD.t231 VDD.n431 146.282
R416 VDD.t158 VDD.n421 146.282
R417 VDD.t312 VDD.n411 146.282
R418 VDD.t249 VDD.n401 146.282
R419 VDD.t36 VDD.n392 146.282
R420 VDD.t195 VDD.n458 144.881
R421 VDD.t34 VDD.n448 144.881
R422 VDD.t452 VDD.n438 144.881
R423 VDD.t74 VDD.n428 144.881
R424 VDD.t48 VDD.n418 144.881
R425 VDD.t164 VDD.n408 144.881
R426 VDD.t492 VDD.n398 144.881
R427 VDD.t340 VDD.n389 144.881
R428 VDD.t233 VDD.n929 143.49
R429 VDD.t270 VDD.n943 143.49
R430 VDD.t193 VDD.n957 143.49
R431 VDD.t387 VDD.n971 143.49
R432 VDD.t154 VDD.n985 143.49
R433 VDD.t383 VDD.n999 143.49
R434 VDD.t434 VDD.n1013 143.49
R435 VDD.n11 VDD.t218 143.49
R436 VDD.n927 VDD.t189 141.511
R437 VDD.n941 VDD.t156 141.511
R438 VDD.n955 VDD.t286 141.511
R439 VDD.n969 VDD.t469 141.511
R440 VDD.n983 VDD.t24 141.511
R441 VDD.n997 VDD.t127 141.511
R442 VDD.n1011 VDD.t82 141.511
R443 VDD.n12 VDD.t28 141.511
R444 VDD.n261 VDD.n256 139.512
R445 VDD.n354 VDD.n77 139.512
R446 VDD.n611 VDD.n606 139.512
R447 VDD.n634 VDD.n557 139.512
R448 VDD.n912 VDD.t288 135.981
R449 VDD.n897 VDD.t258 135.981
R450 VDD.n882 VDD.t496 135.981
R451 VDD.n867 VDD.t413 135.981
R452 VDD.n852 VDD.t338 135.981
R453 VDD.n837 VDD.t292 135.981
R454 VDD.n822 VDD.t94 135.981
R455 VDD.n807 VDD.t282 135.981
R456 VDD.n792 VDD.t310 135.981
R457 VDD.n481 VDD.t356 135.981
R458 VDD.n494 VDD.t306 135.981
R459 VDD.n507 VDD.t176 135.981
R460 VDD.n520 VDD.t100 135.981
R461 VDD.n533 VDD.t187 135.981
R462 VDD.n546 VDD.t375 135.981
R463 VDD.n639 VDD.t30 135.981
R464 VDD.t64 VDD.n913 135.049
R465 VDD.t216 VDD.n898 135.049
R466 VDD.t326 VDD.n883 135.049
R467 VDD.t379 VDD.n868 135.049
R468 VDD.t252 VDD.n853 135.049
R469 VDD.t385 VDD.n838 135.049
R470 VDD.t377 VDD.n823 135.049
R471 VDD.t436 VDD.n808 135.049
R472 VDD.t56 VDD.n793 135.049
R473 VDD.n707 VDD.t262 135.049
R474 VDD.n706 VDD.t334 135.049
R475 VDD.n696 VDD.t133 135.049
R476 VDD.n695 VDD.t237 135.049
R477 VDD.n685 VDD.t465 135.049
R478 VDD.n684 VDD.t212 135.049
R479 VDD.n674 VDD.t460 135.049
R480 VDD.n673 VDD.t318 135.049
R481 VDD.n663 VDD.t244 135.049
R482 VDD.n662 VDD.t431 135.049
R483 VDD.n652 VDD.t119 135.049
R484 VDD.n651 VDD.t32 135.049
R485 VDD.n641 VDD.t467 135.049
R486 VDD.n914 VDD.t268 132.256
R487 VDD.n899 VDD.t442 132.256
R488 VDD.n884 VDD.t129 132.256
R489 VDD.n869 VDD.t346 132.256
R490 VDD.n854 VDD.t500 132.256
R491 VDD.n839 VDD.t125 132.256
R492 VDD.n824 VDD.t448 132.256
R493 VDD.n809 VDD.t183 132.256
R494 VDD.n794 VDD.t117 132.256
R495 VDD.t417 VDD.n482 132.256
R496 VDD.t322 VDD.n495 132.256
R497 VDD.t300 VDD.n508 132.256
R498 VDD.t115 VDD.n521 132.256
R499 VDD.t477 VDD.n534 132.256
R500 VDD.t80 VDD.n547 132.256
R501 VDD.t104 VDD.n640 132.256
R502 VDD.n346 VDD.n87 120.178
R503 VDD.n91 VDD.n89 120.178
R504 VDD.n339 VDD.n94 120.178
R505 VDD.n98 VDD.n96 120.178
R506 VDD.n332 VDD.n101 120.178
R507 VDD.n105 VDD.n103 120.178
R508 VDD.n325 VDD.n108 120.178
R509 VDD.n112 VDD.n110 120.178
R510 VDD.n318 VDD.n115 120.178
R511 VDD.n119 VDD.n117 120.178
R512 VDD.n311 VDD.n122 120.178
R513 VDD.n126 VDD.n124 120.178
R514 VDD.n304 VDD.n129 120.178
R515 VDD.n133 VDD.n131 120.178
R516 VDD.n297 VDD.n136 120.178
R517 VDD.n140 VDD.n138 120.178
R518 VDD.n290 VDD.n143 120.178
R519 VDD.n147 VDD.n145 120.178
R520 VDD.n283 VDD.n150 120.178
R521 VDD.n154 VDD.n152 120.178
R522 VDD.n276 VDD.n157 120.178
R523 VDD.n161 VDD.n159 120.178
R524 VDD.n269 VDD.n164 120.178
R525 VDD.n168 VDD.n166 120.178
R526 VDD.n262 VDD.n171 120.178
R527 VDD.n84 VDD.n82 120.178
R528 VDD.n353 VDD.n80 120.178
R529 VDD.n626 VDD.n567 120.178
R530 VDD.n571 VDD.n569 120.178
R531 VDD.n619 VDD.n574 120.178
R532 VDD.n578 VDD.n576 120.178
R533 VDD.n612 VDD.n581 120.178
R534 VDD.n564 VDD.n562 120.178
R535 VDD.n633 VDD.n560 120.178
R536 VDD VDD.n706 108.04
R537 VDD VDD.n695 108.04
R538 VDD VDD.n684 108.04
R539 VDD VDD.n673 108.04
R540 VDD VDD.n662 108.04
R541 VDD VDD.n651 108.04
R542 VDD.t260 VDD.t296 87.0838
R543 VDD.t180 VDD.t260 87.0838
R544 VDD.t189 VDD.t180 87.0838
R545 VDD.t251 VDD.t233 87.0838
R546 VDD.t290 VDD.t251 87.0838
R547 VDD.t348 VDD.t290 87.0838
R548 VDD.t397 VDD.t342 87.0838
R549 VDD.t494 VDD.t397 87.0838
R550 VDD.t156 VDD.t494 87.0838
R551 VDD.t10 VDD.t270 87.0838
R552 VDD.t225 VDD.t10 87.0838
R553 VDD.t135 VDD.t225 87.0838
R554 VDD.t137 VDD.t444 87.0838
R555 VDD.t248 VDD.t137 87.0838
R556 VDD.t286 VDD.t248 87.0838
R557 VDD.t149 VDD.t193 87.0838
R558 VDD.t458 VDD.t149 87.0838
R559 VDD.t274 VDD.t458 87.0838
R560 VDD.t139 VDD.t0 87.0838
R561 VDD.t224 VDD.t139 87.0838
R562 VDD.t469 VDD.t224 87.0838
R563 VDD.t239 VDD.t387 87.0838
R564 VDD.t4 VDD.t239 87.0838
R565 VDD.t141 VDD.t4 87.0838
R566 VDD.t421 VDD.t419 87.0838
R567 VDD.t491 VDD.t421 87.0838
R568 VDD.t24 VDD.t491 87.0838
R569 VDD.t433 VDD.t154 87.0838
R570 VDD.t425 VDD.t433 87.0838
R571 VDD.t427 VDD.t425 87.0838
R572 VDD.t58 VDD.t328 87.0838
R573 VDD.t462 VDD.t58 87.0838
R574 VDD.t127 VDD.t462 87.0838
R575 VDD.t110 VDD.t383 87.0838
R576 VDD.t391 VDD.t110 87.0838
R577 VDD.t389 VDD.t391 87.0838
R578 VDD.t438 VDD.t362 87.0838
R579 VDD.t15 VDD.t438 87.0838
R580 VDD.t82 VDD.t15 87.0838
R581 VDD.t368 VDD.t434 87.0838
R582 VDD.t360 VDD.t368 87.0838
R583 VDD.t366 VDD.t360 87.0838
R584 VDD.t502 VDD.t86 87.0838
R585 VDD.t495 VDD.t502 87.0838
R586 VDD.t28 VDD.t495 87.0838
R587 VDD.t218 VDD.t197 87.0838
R588 VDD.t197 VDD.t222 87.0838
R589 VDD.t222 VDD.t405 87.0838
R590 VDD.n358 VDD.t196 85.2064
R591 VDD.n362 VDD.t35 85.2064
R592 VDD.n366 VDD.t453 85.2064
R593 VDD.n370 VDD.t75 85.2064
R594 VDD.n374 VDD.t49 85.2064
R595 VDD.n378 VDD.t165 85.2064
R596 VDD.n382 VDD.t493 85.2064
R597 VDD.n386 VDD.t341 85.2064
R598 VDD.n75 VDD.t234 85.0216
R599 VDD.n935 VDD.t190 85.0216
R600 VDD.n67 VDD.t271 85.0216
R601 VDD.n949 VDD.t157 85.0216
R602 VDD.n59 VDD.t194 85.0216
R603 VDD.n963 VDD.t287 85.0216
R604 VDD.n51 VDD.t388 85.0216
R605 VDD.n977 VDD.t470 85.0216
R606 VDD.n43 VDD.t155 85.0216
R607 VDD.n991 VDD.t25 85.0216
R608 VDD.n35 VDD.t384 85.0216
R609 VDD.n1005 VDD.t128 85.0216
R610 VDD.n27 VDD.t435 85.0216
R611 VDD.n1019 VDD.t83 85.0216
R612 VDD.n18 VDD.t219 85.0216
R613 VDD.n3 VDD.t29 85.0216
R614 VDD.n259 VDD.t161 84.7934
R615 VDD.n169 VDD.t408 84.7934
R616 VDD.n266 VDD.t285 84.7934
R617 VDD.n162 VDD.t124 84.7934
R618 VDD.n273 VDD.t241 84.7934
R619 VDD.n155 VDD.t163 84.7934
R620 VDD.n280 VDD.t14 84.7934
R621 VDD.n148 VDD.t53 84.7934
R622 VDD.n287 VDD.t201 84.7934
R623 VDD.n141 VDD.t205 84.7934
R624 VDD.n294 VDD.t199 84.7934
R625 VDD.n134 VDD.t203 84.7934
R626 VDD.n301 VDD.t303 84.7934
R627 VDD.n127 VDD.t107 84.7934
R628 VDD.n308 VDD.t43 84.7934
R629 VDD.n120 VDD.t265 84.7934
R630 VDD.n315 VDD.t89 84.7934
R631 VDD.n113 VDD.t169 84.7934
R632 VDD.n322 VDD.t7 84.7934
R633 VDD.n106 VDD.t109 84.7934
R634 VDD.n329 VDD.t488 84.7934
R635 VDD.n99 VDD.t333 84.7934
R636 VDD.n336 VDD.t167 84.7934
R637 VDD.n92 VDD.t85 84.7934
R638 VDD.n343 VDD.t305 84.7934
R639 VDD.n85 VDD.t267 84.7934
R640 VDD.n350 VDD.t91 84.7934
R641 VDD.n78 VDD.t447 84.7934
R642 VDD.n609 VDD.t192 84.7934
R643 VDD.n579 VDD.t17 84.7934
R644 VDD.n616 VDD.t23 84.7934
R645 VDD.n572 VDD.t21 84.7934
R646 VDD.n623 VDD.t19 84.7934
R647 VDD.n565 VDD.t69 84.7934
R648 VDD.n630 VDD.t277 84.7934
R649 VDD.n558 VDD.t476 84.7934
R650 VDD.n360 VDD.t179 84.7281
R651 VDD.n359 VDD.t209 84.7281
R652 VDD.n358 VDD.t132 84.7281
R653 VDD.n364 VDD.t27 84.7281
R654 VDD.n363 VDD.t396 84.7281
R655 VDD.n362 VDD.t151 84.7281
R656 VDD.n368 VDD.t215 84.7281
R657 VDD.n367 VDD.t484 84.7281
R658 VDD.n366 VDD.t228 84.7281
R659 VDD.n372 VDD.t232 84.7281
R660 VDD.n371 VDD.t144 84.7281
R661 VDD.n370 VDD.t3 84.7281
R662 VDD.n376 VDD.t159 84.7281
R663 VDD.n375 VDD.t430 84.7281
R664 VDD.n374 VDD.t416 84.7281
R665 VDD.n380 VDD.t313 84.7281
R666 VDD.n379 VDD.t455 84.7281
R667 VDD.n378 VDD.t351 84.7281
R668 VDD.n384 VDD.t250 84.7281
R669 VDD.n383 VDD.t230 84.7281
R670 VDD.n382 VDD.t365 84.7281
R671 VDD.n388 VDD.t37 84.7281
R672 VDD.n387 VDD.t39 84.7281
R673 VDD.n386 VDD.t221 84.7281
R674 VDD.t294 VDD.t210 81.9613
R675 VDD.t479 VDD.t294 81.9613
R676 VDD.t288 VDD.t479 81.9613
R677 VDD.t268 VDD.t450 81.9613
R678 VDD.t450 VDD.t8 81.9613
R679 VDD.t8 VDD.t64 81.9613
R680 VDD.t185 VDD.t369 81.9613
R681 VDD.t96 VDD.t185 81.9613
R682 VDD.t258 VDD.t96 81.9613
R683 VDD.t442 VDD.t98 81.9613
R684 VDD.t98 VDD.t254 81.9613
R685 VDD.t254 VDD.t216 81.9613
R686 VDD.t76 VDD.t181 81.9613
R687 VDD.t78 VDD.t76 81.9613
R688 VDD.t496 VDD.t78 81.9613
R689 VDD.t129 VDD.t354 81.9613
R690 VDD.t354 VDD.t324 81.9613
R691 VDD.t324 VDD.t326 81.9613
R692 VDD.t411 VDD.t481 81.9613
R693 VDD.t358 VDD.t411 81.9613
R694 VDD.t413 VDD.t358 81.9613
R695 VDD.t346 VDD.t11 81.9613
R696 VDD.t11 VDD.t381 81.9613
R697 VDD.t381 VDD.t379 81.9613
R698 VDD.t371 VDD.t473 81.9613
R699 VDD.t463 VDD.t371 81.9613
R700 VDD.t338 VDD.t463 81.9613
R701 VDD.t500 VDD.t399 81.9613
R702 VDD.t399 VDD.t498 81.9613
R703 VDD.t498 VDD.t252 81.9613
R704 VDD.t111 VDD.t298 81.9613
R705 VDD.t330 VDD.t111 81.9613
R706 VDD.t292 VDD.t330 81.9613
R707 VDD.t125 VDD.t256 81.9613
R708 VDD.t256 VDD.t54 81.9613
R709 VDD.t54 VDD.t385 81.9613
R710 VDD.t62 VDD.t92 81.9613
R711 VDD.t121 VDD.t62 81.9613
R712 VDD.t94 VDD.t121 81.9613
R713 VDD.t448 VDD.t172 81.9613
R714 VDD.t172 VDD.t46 81.9613
R715 VDD.t46 VDD.t377 81.9613
R716 VDD.t70 VDD.t280 81.9613
R717 VDD.t278 VDD.t70 81.9613
R718 VDD.t282 VDD.t278 81.9613
R719 VDD.t183 VDD.t235 81.9613
R720 VDD.t235 VDD.t336 81.9613
R721 VDD.t336 VDD.t436 81.9613
R722 VDD.t393 VDD.t409 81.9613
R723 VDD.t308 VDD.t393 81.9613
R724 VDD.t310 VDD.t308 81.9613
R725 VDD.t117 VDD.t489 81.9613
R726 VDD.t489 VDD.t72 81.9613
R727 VDD.t72 VDD.t56 81.9613
R728 VDD.t145 VDD.t403 81.9613
R729 VDD.t403 VDD.t320 81.9613
R730 VDD.t320 VDD.t356 81.9613
R731 VDD.t344 VDD.t417 81.9613
R732 VDD.t423 VDD.t344 81.9613
R733 VDD.t262 VDD.t423 81.9613
R734 VDD.t471 VDD.t334 81.9613
R735 VDD.t206 VDD.t471 81.9613
R736 VDD.t306 VDD.t206 81.9613
R737 VDD.t147 VDD.t322 81.9613
R738 VDD.t401 VDD.t147 81.9613
R739 VDD.t133 VDD.t401 81.9613
R740 VDD.t50 VDD.t237 81.9613
R741 VDD.t174 VDD.t50 81.9613
R742 VDD.t176 VDD.t174 81.9613
R743 VDD.t242 VDD.t300 81.9613
R744 VDD.t102 VDD.t242 81.9613
R745 VDD.t465 VDD.t102 81.9613
R746 VDD.t66 VDD.t212 81.9613
R747 VDD.t314 VDD.t66 81.9613
R748 VDD.t100 VDD.t314 81.9613
R749 VDD.t44 VDD.t115 81.9613
R750 VDD.t352 VDD.t44 81.9613
R751 VDD.t460 VDD.t352 81.9613
R752 VDD.t113 VDD.t318 81.9613
R753 VDD.t456 VDD.t113 81.9613
R754 VDD.t187 VDD.t456 81.9613
R755 VDD.t316 VDD.t477 81.9613
R756 VDD.t272 VDD.t316 81.9613
R757 VDD.t244 VDD.t272 81.9613
R758 VDD.t373 VDD.t431 81.9613
R759 VDD.t60 VDD.t373 81.9613
R760 VDD.t375 VDD.t60 81.9613
R761 VDD.t170 VDD.t80 81.9613
R762 VDD.t152 VDD.t170 81.9613
R763 VDD.t119 VDD.t152 81.9613
R764 VDD.t440 VDD.t32 81.9613
R765 VDD.t246 VDD.t440 81.9613
R766 VDD.t30 VDD.t246 81.9613
R767 VDD.t40 VDD.t104 81.9613
R768 VDD.t485 VDD.t40 81.9613
R769 VDD.t467 VDD.t485 81.9613
R770 VDD.t131 VDD.t195 78.5719
R771 VDD.t208 VDD.t178 78.5719
R772 VDD.t150 VDD.t34 78.5719
R773 VDD.t395 VDD.t26 78.5719
R774 VDD.t227 VDD.t452 78.5719
R775 VDD.t483 VDD.t214 78.5719
R776 VDD.t2 VDD.t74 78.5719
R777 VDD.t143 VDD.t231 78.5719
R778 VDD.t415 VDD.t48 78.5719
R779 VDD.t429 VDD.t158 78.5719
R780 VDD.t350 VDD.t164 78.5719
R781 VDD.t454 VDD.t312 78.5719
R782 VDD.t364 VDD.t492 78.5719
R783 VDD.t229 VDD.t249 78.5719
R784 VDD.t220 VDD.t340 78.5719
R785 VDD.t38 VDD.t36 78.5719
R786 VDD.n919 VDD.n716 75.7173
R787 VDD.n918 VDD.n717 75.7173
R788 VDD.n719 VDD.n718 75.7173
R789 VDD.n907 VDD.n906 75.7173
R790 VDD.n904 VDD.n724 75.7173
R791 VDD.n903 VDD.n725 75.7173
R792 VDD.n727 VDD.n726 75.7173
R793 VDD.n892 VDD.n891 75.7173
R794 VDD.n889 VDD.n732 75.7173
R795 VDD.n888 VDD.n733 75.7173
R796 VDD.n735 VDD.n734 75.7173
R797 VDD.n877 VDD.n876 75.7173
R798 VDD.n874 VDD.n740 75.7173
R799 VDD.n873 VDD.n741 75.7173
R800 VDD.n743 VDD.n742 75.7173
R801 VDD.n862 VDD.n861 75.7173
R802 VDD.n859 VDD.n748 75.7173
R803 VDD.n858 VDD.n749 75.7173
R804 VDD.n751 VDD.n750 75.7173
R805 VDD.n847 VDD.n846 75.7173
R806 VDD.n844 VDD.n756 75.7173
R807 VDD.n843 VDD.n757 75.7173
R808 VDD.n759 VDD.n758 75.7173
R809 VDD.n832 VDD.n831 75.7173
R810 VDD.n829 VDD.n764 75.7173
R811 VDD.n828 VDD.n765 75.7173
R812 VDD.n767 VDD.n766 75.7173
R813 VDD.n817 VDD.n816 75.7173
R814 VDD.n814 VDD.n772 75.7173
R815 VDD.n813 VDD.n773 75.7173
R816 VDD.n775 VDD.n774 75.7173
R817 VDD.n802 VDD.n801 75.7173
R818 VDD.n799 VDD.n780 75.7173
R819 VDD.n798 VDD.n781 75.7173
R820 VDD.n783 VDD.n782 75.7173
R821 VDD.n788 VDD.n787 75.7173
R822 VDD.n556 VDD.n555 75.7173
R823 VDD.n553 VDD.n552 75.7173
R824 VDD.n646 VDD.n551 75.7173
R825 VDD.n647 VDD.n550 75.7173
R826 VDD.n543 VDD.n542 75.7173
R827 VDD.n540 VDD.n539 75.7173
R828 VDD.n657 VDD.n538 75.7173
R829 VDD.n658 VDD.n537 75.7173
R830 VDD.n530 VDD.n529 75.7173
R831 VDD.n527 VDD.n526 75.7173
R832 VDD.n668 VDD.n525 75.7173
R833 VDD.n669 VDD.n524 75.7173
R834 VDD.n517 VDD.n516 75.7173
R835 VDD.n514 VDD.n513 75.7173
R836 VDD.n679 VDD.n512 75.7173
R837 VDD.n680 VDD.n511 75.7173
R838 VDD.n504 VDD.n503 75.7173
R839 VDD.n501 VDD.n500 75.7173
R840 VDD.n690 VDD.n499 75.7173
R841 VDD.n691 VDD.n498 75.7173
R842 VDD.n491 VDD.n490 75.7173
R843 VDD.n488 VDD.n487 75.7173
R844 VDD.n701 VDD.n486 75.7173
R845 VDD.n702 VDD.n485 75.7173
R846 VDD.n476 VDD.n475 75.7173
R847 VDD.n472 VDD.n471 75.7173
R848 VDD.n712 VDD.n470 75.7173
R849 VDD.n713 VDD.n469 75.7173
R850 VDD.n76 VDD.n74 75.5
R851 VDD.n936 VDD.n70 75.5
R852 VDD.n68 VDD.n66 75.5
R853 VDD.n950 VDD.n62 75.5
R854 VDD.n60 VDD.n58 75.5
R855 VDD.n964 VDD.n54 75.5
R856 VDD.n52 VDD.n50 75.5
R857 VDD.n978 VDD.n46 75.5
R858 VDD.n44 VDD.n42 75.5
R859 VDD.n992 VDD.n38 75.5
R860 VDD.n36 VDD.n34 75.5
R861 VDD.n1006 VDD.n30 75.5
R862 VDD.n28 VDD.n26 75.5
R863 VDD.n1020 VDD.n22 75.5
R864 VDD.n19 VDD.n1 75.5
R865 VDD.n5 VDD.n4 75.5
R866 VDD.n913 VDD 50.2946
R867 VDD.n898 VDD 50.2946
R868 VDD.n883 VDD 50.2946
R869 VDD.n868 VDD 50.2946
R870 VDD.n853 VDD 50.2946
R871 VDD.n838 VDD 50.2946
R872 VDD.n823 VDD 50.2946
R873 VDD.n808 VDD 50.2946
R874 VDD.n793 VDD 50.2946
R875 VDD.n707 VDD 50.2946
R876 VDD.n696 VDD 50.2946
R877 VDD.n685 VDD 50.2946
R878 VDD.n674 VDD 50.2946
R879 VDD.n663 VDD 50.2946
R880 VDD.n652 VDD 50.2946
R881 VDD.n641 VDD 50.2946
R882 VDD.n354 VDD.n79 46.2505
R883 VDD.n352 VDD.n81 46.2505
R884 VDD.t90 VDD.n81 46.2505
R885 VDD.n347 VDD.n86 46.2505
R886 VDD.t266 VDD.n86 46.2505
R887 VDD.n345 VDD.n88 46.2505
R888 VDD.t304 VDD.n88 46.2505
R889 VDD.n340 VDD.n93 46.2505
R890 VDD.t84 VDD.n93 46.2505
R891 VDD.n338 VDD.n95 46.2505
R892 VDD.t166 VDD.n95 46.2505
R893 VDD.n333 VDD.n100 46.2505
R894 VDD.t332 VDD.n100 46.2505
R895 VDD.n331 VDD.n102 46.2505
R896 VDD.t487 VDD.n102 46.2505
R897 VDD.n326 VDD.n107 46.2505
R898 VDD.t108 VDD.n107 46.2505
R899 VDD.n324 VDD.n109 46.2505
R900 VDD.t6 VDD.n109 46.2505
R901 VDD.n319 VDD.n114 46.2505
R902 VDD.t168 VDD.n114 46.2505
R903 VDD.n317 VDD.n116 46.2505
R904 VDD.t88 VDD.n116 46.2505
R905 VDD.n312 VDD.n121 46.2505
R906 VDD.t264 VDD.n121 46.2505
R907 VDD.n310 VDD.n123 46.2505
R908 VDD.t42 VDD.n123 46.2505
R909 VDD.n305 VDD.n128 46.2505
R910 VDD.t106 VDD.n128 46.2505
R911 VDD.n303 VDD.n130 46.2505
R912 VDD.t302 VDD.n130 46.2505
R913 VDD.n298 VDD.n135 46.2505
R914 VDD.t202 VDD.n135 46.2505
R915 VDD.n296 VDD.n137 46.2505
R916 VDD.t198 VDD.n137 46.2505
R917 VDD.n291 VDD.n142 46.2505
R918 VDD.t204 VDD.n142 46.2505
R919 VDD.n289 VDD.n144 46.2505
R920 VDD.t200 VDD.n144 46.2505
R921 VDD.n284 VDD.n149 46.2505
R922 VDD.t52 VDD.n149 46.2505
R923 VDD.n282 VDD.n151 46.2505
R924 VDD.t13 VDD.n151 46.2505
R925 VDD.n277 VDD.n156 46.2505
R926 VDD.t162 VDD.n156 46.2505
R927 VDD.n275 VDD.n158 46.2505
R928 VDD.t240 VDD.n158 46.2505
R929 VDD.n270 VDD.n163 46.2505
R930 VDD.t123 VDD.n163 46.2505
R931 VDD.n268 VDD.n165 46.2505
R932 VDD.t284 VDD.n165 46.2505
R933 VDD.n263 VDD.n170 46.2505
R934 VDD.t407 VDD.n170 46.2505
R935 VDD.n261 VDD.n172 46.2505
R936 VDD.n634 VDD.n559 46.2505
R937 VDD.n632 VDD.n561 46.2505
R938 VDD.t276 VDD.n561 46.2505
R939 VDD.n627 VDD.n566 46.2505
R940 VDD.t68 VDD.n566 46.2505
R941 VDD.n625 VDD.n568 46.2505
R942 VDD.t18 VDD.n568 46.2505
R943 VDD.n620 VDD.n573 46.2505
R944 VDD.t20 VDD.n573 46.2505
R945 VDD.n618 VDD.n575 46.2505
R946 VDD.t22 VDD.n575 46.2505
R947 VDD.n613 VDD.n580 46.2505
R948 VDD.t16 VDD.n580 46.2505
R949 VDD.n611 VDD.n582 46.2505
R950 VDD.n173 VDD.n79 39.3924
R951 VDD.n255 VDD.n172 39.3924
R952 VDD.n583 VDD.n559 39.3924
R953 VDD.n605 VDD.n582 39.3924
R954 VDD.n463 VDD.n462 38.0519
R955 VDD.n453 VDD.n452 38.0519
R956 VDD.n443 VDD.n442 38.0519
R957 VDD.n433 VDD.n432 38.0519
R958 VDD.n423 VDD.n422 38.0519
R959 VDD.n413 VDD.n412 38.0519
R960 VDD.n403 VDD.n402 38.0519
R961 VDD.n394 VDD.n393 38.0519
R962 VDD.n253 VDD.n171 20.5561
R963 VDD.n254 VDD.n253 20.5561
R964 VDD.n250 VDD.n168 20.5561
R965 VDD.n251 VDD.n250 20.5561
R966 VDD.n247 VDD.n164 20.5561
R967 VDD.n248 VDD.n247 20.5561
R968 VDD.n244 VDD.n161 20.5561
R969 VDD.n245 VDD.n244 20.5561
R970 VDD.n241 VDD.n157 20.5561
R971 VDD.n242 VDD.n241 20.5561
R972 VDD.n238 VDD.n154 20.5561
R973 VDD.n239 VDD.n238 20.5561
R974 VDD.n235 VDD.n150 20.5561
R975 VDD.n236 VDD.n235 20.5561
R976 VDD.n232 VDD.n147 20.5561
R977 VDD.n233 VDD.n232 20.5561
R978 VDD.n229 VDD.n143 20.5561
R979 VDD.n230 VDD.n229 20.5561
R980 VDD.n226 VDD.n140 20.5561
R981 VDD.n227 VDD.n226 20.5561
R982 VDD.n223 VDD.n136 20.5561
R983 VDD.n224 VDD.n223 20.5561
R984 VDD.n220 VDD.n133 20.5561
R985 VDD.n221 VDD.n220 20.5561
R986 VDD.n217 VDD.n129 20.5561
R987 VDD.n218 VDD.n217 20.5561
R988 VDD.n214 VDD.n126 20.5561
R989 VDD.n215 VDD.n214 20.5561
R990 VDD.n211 VDD.n122 20.5561
R991 VDD.n212 VDD.n211 20.5561
R992 VDD.n208 VDD.n119 20.5561
R993 VDD.n209 VDD.n208 20.5561
R994 VDD.n205 VDD.n115 20.5561
R995 VDD.n206 VDD.n205 20.5561
R996 VDD.n202 VDD.n112 20.5561
R997 VDD.n203 VDD.n202 20.5561
R998 VDD.n199 VDD.n108 20.5561
R999 VDD.n200 VDD.n199 20.5561
R1000 VDD.n196 VDD.n105 20.5561
R1001 VDD.n197 VDD.n196 20.5561
R1002 VDD.n193 VDD.n101 20.5561
R1003 VDD.n194 VDD.n193 20.5561
R1004 VDD.n190 VDD.n98 20.5561
R1005 VDD.n191 VDD.n190 20.5561
R1006 VDD.n187 VDD.n94 20.5561
R1007 VDD.n188 VDD.n187 20.5561
R1008 VDD.n184 VDD.n91 20.5561
R1009 VDD.n185 VDD.n184 20.5561
R1010 VDD.n181 VDD.n87 20.5561
R1011 VDD.n182 VDD.n181 20.5561
R1012 VDD.n178 VDD.n84 20.5561
R1013 VDD.n179 VDD.n178 20.5561
R1014 VDD.n175 VDD.n80 20.5561
R1015 VDD.n176 VDD.n175 20.5561
R1016 VDD.n603 VDD.n581 20.5561
R1017 VDD.n604 VDD.n603 20.5561
R1018 VDD.n600 VDD.n578 20.5561
R1019 VDD.n601 VDD.n600 20.5561
R1020 VDD.n597 VDD.n574 20.5561
R1021 VDD.n598 VDD.n597 20.5561
R1022 VDD.n594 VDD.n571 20.5561
R1023 VDD.n595 VDD.n594 20.5561
R1024 VDD.n591 VDD.n567 20.5561
R1025 VDD.n592 VDD.n591 20.5561
R1026 VDD.n588 VDD.n564 20.5561
R1027 VDD.n589 VDD.n588 20.5561
R1028 VDD.n585 VDD.n560 20.5561
R1029 VDD.n586 VDD.n585 20.5561
R1030 VDD.n931 VDD.n930 20.5561
R1031 VDD.n928 VDD.n73 20.5561
R1032 VDD.n929 VDD.n928 20.5561
R1033 VDD.n926 VDD.n69 20.5561
R1034 VDD.n945 VDD.n944 20.5561
R1035 VDD.n942 VDD.n65 20.5561
R1036 VDD.n943 VDD.n942 20.5561
R1037 VDD.n940 VDD.n61 20.5561
R1038 VDD.n959 VDD.n958 20.5561
R1039 VDD.n956 VDD.n57 20.5561
R1040 VDD.n957 VDD.n956 20.5561
R1041 VDD.n954 VDD.n53 20.5561
R1042 VDD.n973 VDD.n972 20.5561
R1043 VDD.n970 VDD.n49 20.5561
R1044 VDD.n971 VDD.n970 20.5561
R1045 VDD.n968 VDD.n45 20.5561
R1046 VDD.n987 VDD.n986 20.5561
R1047 VDD.n984 VDD.n41 20.5561
R1048 VDD.n985 VDD.n984 20.5561
R1049 VDD.n982 VDD.n37 20.5561
R1050 VDD.n1001 VDD.n1000 20.5561
R1051 VDD.n998 VDD.n33 20.5561
R1052 VDD.n999 VDD.n998 20.5561
R1053 VDD.n996 VDD.n29 20.5561
R1054 VDD.n1015 VDD.n1014 20.5561
R1055 VDD.n1012 VDD.n25 20.5561
R1056 VDD.n1013 VDD.n1012 20.5561
R1057 VDD.n1010 VDD.n21 20.5561
R1058 VDD.n9 VDD.n0 20.5561
R1059 VDD.n10 VDD.n2 20.5561
R1060 VDD.n11 VDD.n10 20.5561
R1061 VDD.n7 VDD.n6 20.5561
R1062 VDD.n354 VDD.n353 19.3338
R1063 VDD.n353 VDD.n352 19.3338
R1064 VDD.n352 VDD.n82 19.3338
R1065 VDD.n347 VDD.n82 19.3338
R1066 VDD.n347 VDD.n346 19.3338
R1067 VDD.n346 VDD.n345 19.3338
R1068 VDD.n345 VDD.n89 19.3338
R1069 VDD.n340 VDD.n89 19.3338
R1070 VDD.n340 VDD.n339 19.3338
R1071 VDD.n339 VDD.n338 19.3338
R1072 VDD.n338 VDD.n96 19.3338
R1073 VDD.n333 VDD.n96 19.3338
R1074 VDD.n333 VDD.n332 19.3338
R1075 VDD.n332 VDD.n331 19.3338
R1076 VDD.n331 VDD.n103 19.3338
R1077 VDD.n326 VDD.n103 19.3338
R1078 VDD.n326 VDD.n325 19.3338
R1079 VDD.n325 VDD.n324 19.3338
R1080 VDD.n324 VDD.n110 19.3338
R1081 VDD.n319 VDD.n110 19.3338
R1082 VDD.n319 VDD.n318 19.3338
R1083 VDD.n318 VDD.n317 19.3338
R1084 VDD.n317 VDD.n117 19.3338
R1085 VDD.n312 VDD.n117 19.3338
R1086 VDD.n312 VDD.n311 19.3338
R1087 VDD.n311 VDD.n310 19.3338
R1088 VDD.n310 VDD.n124 19.3338
R1089 VDD.n305 VDD.n124 19.3338
R1090 VDD.n305 VDD.n304 19.3338
R1091 VDD.n304 VDD.n303 19.3338
R1092 VDD.n303 VDD.n131 19.3338
R1093 VDD.n298 VDD.n131 19.3338
R1094 VDD.n298 VDD.n297 19.3338
R1095 VDD.n297 VDD.n296 19.3338
R1096 VDD.n296 VDD.n138 19.3338
R1097 VDD.n291 VDD.n138 19.3338
R1098 VDD.n291 VDD.n290 19.3338
R1099 VDD.n290 VDD.n289 19.3338
R1100 VDD.n289 VDD.n145 19.3338
R1101 VDD.n284 VDD.n145 19.3338
R1102 VDD.n284 VDD.n283 19.3338
R1103 VDD.n283 VDD.n282 19.3338
R1104 VDD.n282 VDD.n152 19.3338
R1105 VDD.n277 VDD.n152 19.3338
R1106 VDD.n277 VDD.n276 19.3338
R1107 VDD.n276 VDD.n275 19.3338
R1108 VDD.n275 VDD.n159 19.3338
R1109 VDD.n270 VDD.n159 19.3338
R1110 VDD.n270 VDD.n269 19.3338
R1111 VDD.n269 VDD.n268 19.3338
R1112 VDD.n268 VDD.n166 19.3338
R1113 VDD.n263 VDD.n166 19.3338
R1114 VDD.n263 VDD.n262 19.3338
R1115 VDD.n262 VDD.n261 19.3338
R1116 VDD.n634 VDD.n633 19.3338
R1117 VDD.n633 VDD.n632 19.3338
R1118 VDD.n632 VDD.n562 19.3338
R1119 VDD.n627 VDD.n562 19.3338
R1120 VDD.n627 VDD.n626 19.3338
R1121 VDD.n626 VDD.n625 19.3338
R1122 VDD.n625 VDD.n569 19.3338
R1123 VDD.n620 VDD.n569 19.3338
R1124 VDD.n620 VDD.n619 19.3338
R1125 VDD.n619 VDD.n618 19.3338
R1126 VDD.n618 VDD.n576 19.3338
R1127 VDD.n613 VDD.n576 19.3338
R1128 VDD.n613 VDD.n612 19.3338
R1129 VDD.n612 VDD.n611 19.3338
R1130 VDD.n722 VDD.n715 16.8187
R1131 VDD.n913 VDD.n722 16.8187
R1132 VDD.n912 VDD.n911 16.8187
R1133 VDD.n910 VDD.n909 16.8187
R1134 VDD.n730 VDD.n723 16.8187
R1135 VDD.n898 VDD.n730 16.8187
R1136 VDD.n897 VDD.n896 16.8187
R1137 VDD.n895 VDD.n894 16.8187
R1138 VDD.n738 VDD.n731 16.8187
R1139 VDD.n883 VDD.n738 16.8187
R1140 VDD.n882 VDD.n881 16.8187
R1141 VDD.n880 VDD.n879 16.8187
R1142 VDD.n746 VDD.n739 16.8187
R1143 VDD.n868 VDD.n746 16.8187
R1144 VDD.n867 VDD.n866 16.8187
R1145 VDD.n865 VDD.n864 16.8187
R1146 VDD.n754 VDD.n747 16.8187
R1147 VDD.n853 VDD.n754 16.8187
R1148 VDD.n852 VDD.n851 16.8187
R1149 VDD.n850 VDD.n849 16.8187
R1150 VDD.n762 VDD.n755 16.8187
R1151 VDD.n838 VDD.n762 16.8187
R1152 VDD.n837 VDD.n836 16.8187
R1153 VDD.n835 VDD.n834 16.8187
R1154 VDD.n770 VDD.n763 16.8187
R1155 VDD.n823 VDD.n770 16.8187
R1156 VDD.n822 VDD.n821 16.8187
R1157 VDD.n820 VDD.n819 16.8187
R1158 VDD.n778 VDD.n771 16.8187
R1159 VDD.n808 VDD.n778 16.8187
R1160 VDD.n807 VDD.n806 16.8187
R1161 VDD.n805 VDD.n804 16.8187
R1162 VDD.n786 VDD.n779 16.8187
R1163 VDD.n793 VDD.n786 16.8187
R1164 VDD.n792 VDD.n791 16.8187
R1165 VDD.n790 VDD.n789 16.8187
R1166 VDD.n698 VDD.n697 16.8187
R1167 VDD.n697 VDD.n696 16.8187
R1168 VDD.n494 VDD.n493 16.8187
R1169 VDD.n705 VDD.n704 16.8187
R1170 VDD.n706 VDD.n705 16.8187
R1171 VDD.n687 VDD.n686 16.8187
R1172 VDD.n686 VDD.n685 16.8187
R1173 VDD.n507 VDD.n506 16.8187
R1174 VDD.n694 VDD.n693 16.8187
R1175 VDD.n695 VDD.n694 16.8187
R1176 VDD.n676 VDD.n675 16.8187
R1177 VDD.n675 VDD.n674 16.8187
R1178 VDD.n520 VDD.n519 16.8187
R1179 VDD.n683 VDD.n682 16.8187
R1180 VDD.n684 VDD.n683 16.8187
R1181 VDD.n665 VDD.n664 16.8187
R1182 VDD.n664 VDD.n663 16.8187
R1183 VDD.n533 VDD.n532 16.8187
R1184 VDD.n672 VDD.n671 16.8187
R1185 VDD.n673 VDD.n672 16.8187
R1186 VDD.n654 VDD.n653 16.8187
R1187 VDD.n653 VDD.n652 16.8187
R1188 VDD.n546 VDD.n545 16.8187
R1189 VDD.n661 VDD.n660 16.8187
R1190 VDD.n662 VDD.n661 16.8187
R1191 VDD.n643 VDD.n642 16.8187
R1192 VDD.n642 VDD.n641 16.8187
R1193 VDD.n639 VDD.n638 16.8187
R1194 VDD.n650 VDD.n649 16.8187
R1195 VDD.n651 VDD.n650 16.8187
R1196 VDD.n709 VDD.n708 16.8187
R1197 VDD.n708 VDD.n707 16.8187
R1198 VDD.n481 VDD.n480 16.8187
R1199 VDD.n478 VDD.n468 16.8187
R1200 VDD.n461 VDD.n357 16.8187
R1201 VDD.n451 VDD.n361 16.8187
R1202 VDD.n441 VDD.n365 16.8187
R1203 VDD.n431 VDD.n369 16.8187
R1204 VDD.n421 VDD.n373 16.8187
R1205 VDD.n411 VDD.n377 16.8187
R1206 VDD.n401 VDD.n381 16.8187
R1207 VDD.n392 VDD.n385 16.8187
R1208 VDD.n462 VDD.n460 12.5005
R1209 VDD.n452 VDD.n450 12.5005
R1210 VDD.n442 VDD.n440 12.5005
R1211 VDD.n432 VDD.n430 12.5005
R1212 VDD.n422 VDD.n420 12.5005
R1213 VDD.n412 VDD.n410 12.5005
R1214 VDD.n402 VDD.n400 12.5005
R1215 VDD.n393 VDD.n391 12.5005
R1216 VDD.n916 VDD.n915 11.563
R1217 VDD.n915 VDD.n914 11.563
R1218 VDD.n901 VDD.n900 11.563
R1219 VDD.n900 VDD.n899 11.563
R1220 VDD.n886 VDD.n885 11.563
R1221 VDD.n885 VDD.n884 11.563
R1222 VDD.n871 VDD.n870 11.563
R1223 VDD.n870 VDD.n869 11.563
R1224 VDD.n856 VDD.n855 11.563
R1225 VDD.n855 VDD.n854 11.563
R1226 VDD.n841 VDD.n840 11.563
R1227 VDD.n840 VDD.n839 11.563
R1228 VDD.n826 VDD.n825 11.563
R1229 VDD.n825 VDD.n824 11.563
R1230 VDD.n811 VDD.n810 11.563
R1231 VDD.n810 VDD.n809 11.563
R1232 VDD.n796 VDD.n795 11.563
R1233 VDD.n795 VDD.n794 11.563
R1234 VDD.n699 VDD.n489 11.563
R1235 VDD.n495 VDD.n489 11.563
R1236 VDD.n688 VDD.n502 11.563
R1237 VDD.n508 VDD.n502 11.563
R1238 VDD.n677 VDD.n515 11.563
R1239 VDD.n521 VDD.n515 11.563
R1240 VDD.n666 VDD.n528 11.563
R1241 VDD.n534 VDD.n528 11.563
R1242 VDD.n655 VDD.n541 11.563
R1243 VDD.n547 VDD.n541 11.563
R1244 VDD.n644 VDD.n554 11.563
R1245 VDD.n640 VDD.n554 11.563
R1246 VDD.n710 VDD.n474 11.563
R1247 VDD.n482 VDD.n474 11.563
R1248 VDD.n716 VDD.t9 9.52217
R1249 VDD.n716 VDD.t65 9.52217
R1250 VDD.n717 VDD.t269 9.52217
R1251 VDD.n717 VDD.t451 9.52217
R1252 VDD.n718 VDD.t480 9.52217
R1253 VDD.n718 VDD.t289 9.52217
R1254 VDD.n906 VDD.t211 9.52217
R1255 VDD.n906 VDD.t295 9.52217
R1256 VDD.n724 VDD.t255 9.52217
R1257 VDD.n724 VDD.t217 9.52217
R1258 VDD.n725 VDD.t443 9.52217
R1259 VDD.n725 VDD.t99 9.52217
R1260 VDD.n726 VDD.t97 9.52217
R1261 VDD.n726 VDD.t259 9.52217
R1262 VDD.n891 VDD.t370 9.52217
R1263 VDD.n891 VDD.t186 9.52217
R1264 VDD.n732 VDD.t325 9.52217
R1265 VDD.n732 VDD.t327 9.52217
R1266 VDD.n733 VDD.t130 9.52217
R1267 VDD.n733 VDD.t355 9.52217
R1268 VDD.n734 VDD.t79 9.52217
R1269 VDD.n734 VDD.t497 9.52217
R1270 VDD.n876 VDD.t182 9.52217
R1271 VDD.n876 VDD.t77 9.52217
R1272 VDD.n740 VDD.t382 9.52217
R1273 VDD.n740 VDD.t380 9.52217
R1274 VDD.n741 VDD.t347 9.52217
R1275 VDD.n741 VDD.t12 9.52217
R1276 VDD.n742 VDD.t359 9.52217
R1277 VDD.n742 VDD.t414 9.52217
R1278 VDD.n861 VDD.t482 9.52217
R1279 VDD.n861 VDD.t412 9.52217
R1280 VDD.n748 VDD.t499 9.52217
R1281 VDD.n748 VDD.t253 9.52217
R1282 VDD.n749 VDD.t501 9.52217
R1283 VDD.n749 VDD.t400 9.52217
R1284 VDD.n750 VDD.t464 9.52217
R1285 VDD.n750 VDD.t339 9.52217
R1286 VDD.n846 VDD.t474 9.52217
R1287 VDD.n846 VDD.t372 9.52217
R1288 VDD.n756 VDD.t55 9.52217
R1289 VDD.n756 VDD.t386 9.52217
R1290 VDD.n757 VDD.t126 9.52217
R1291 VDD.n757 VDD.t257 9.52217
R1292 VDD.n758 VDD.t331 9.52217
R1293 VDD.n758 VDD.t293 9.52217
R1294 VDD.n831 VDD.t299 9.52217
R1295 VDD.n831 VDD.t112 9.52217
R1296 VDD.n764 VDD.t47 9.52217
R1297 VDD.n764 VDD.t378 9.52217
R1298 VDD.n765 VDD.t449 9.52217
R1299 VDD.n765 VDD.t173 9.52217
R1300 VDD.n766 VDD.t122 9.52217
R1301 VDD.n766 VDD.t95 9.52217
R1302 VDD.n816 VDD.t93 9.52217
R1303 VDD.n816 VDD.t63 9.52217
R1304 VDD.n772 VDD.t337 9.52217
R1305 VDD.n772 VDD.t437 9.52217
R1306 VDD.n773 VDD.t184 9.52217
R1307 VDD.n773 VDD.t236 9.52217
R1308 VDD.n774 VDD.t279 9.52217
R1309 VDD.n774 VDD.t283 9.52217
R1310 VDD.n801 VDD.t281 9.52217
R1311 VDD.n801 VDD.t71 9.52217
R1312 VDD.n780 VDD.t73 9.52217
R1313 VDD.n780 VDD.t57 9.52217
R1314 VDD.n781 VDD.t118 9.52217
R1315 VDD.n781 VDD.t490 9.52217
R1316 VDD.n782 VDD.t309 9.52217
R1317 VDD.n782 VDD.t311 9.52217
R1318 VDD.n787 VDD.t410 9.52217
R1319 VDD.n787 VDD.t394 9.52217
R1320 VDD.n555 VDD.t486 9.52217
R1321 VDD.n555 VDD.t468 9.52217
R1322 VDD.n552 VDD.t105 9.52217
R1323 VDD.n552 VDD.t41 9.52217
R1324 VDD.n551 VDD.t247 9.52217
R1325 VDD.n551 VDD.t31 9.52217
R1326 VDD.n550 VDD.t33 9.52217
R1327 VDD.n550 VDD.t441 9.52217
R1328 VDD.n542 VDD.t153 9.52217
R1329 VDD.n542 VDD.t120 9.52217
R1330 VDD.n539 VDD.t81 9.52217
R1331 VDD.n539 VDD.t171 9.52217
R1332 VDD.n538 VDD.t61 9.52217
R1333 VDD.n538 VDD.t376 9.52217
R1334 VDD.n537 VDD.t432 9.52217
R1335 VDD.n537 VDD.t374 9.52217
R1336 VDD.n529 VDD.t273 9.52217
R1337 VDD.n529 VDD.t245 9.52217
R1338 VDD.n526 VDD.t478 9.52217
R1339 VDD.n526 VDD.t317 9.52217
R1340 VDD.n525 VDD.t457 9.52217
R1341 VDD.n525 VDD.t188 9.52217
R1342 VDD.n524 VDD.t319 9.52217
R1343 VDD.n524 VDD.t114 9.52217
R1344 VDD.n516 VDD.t353 9.52217
R1345 VDD.n516 VDD.t461 9.52217
R1346 VDD.n513 VDD.t116 9.52217
R1347 VDD.n513 VDD.t45 9.52217
R1348 VDD.n512 VDD.t315 9.52217
R1349 VDD.n512 VDD.t101 9.52217
R1350 VDD.n511 VDD.t213 9.52217
R1351 VDD.n511 VDD.t67 9.52217
R1352 VDD.n503 VDD.t103 9.52217
R1353 VDD.n503 VDD.t466 9.52217
R1354 VDD.n500 VDD.t301 9.52217
R1355 VDD.n500 VDD.t243 9.52217
R1356 VDD.n499 VDD.t175 9.52217
R1357 VDD.n499 VDD.t177 9.52217
R1358 VDD.n498 VDD.t238 9.52217
R1359 VDD.n498 VDD.t51 9.52217
R1360 VDD.n490 VDD.t402 9.52217
R1361 VDD.n490 VDD.t134 9.52217
R1362 VDD.n487 VDD.t323 9.52217
R1363 VDD.n487 VDD.t148 9.52217
R1364 VDD.n486 VDD.t207 9.52217
R1365 VDD.n486 VDD.t307 9.52217
R1366 VDD.n485 VDD.t335 9.52217
R1367 VDD.n485 VDD.t472 9.52217
R1368 VDD.n475 VDD.t424 9.52217
R1369 VDD.n475 VDD.t263 9.52217
R1370 VDD.n471 VDD.t418 9.52217
R1371 VDD.n471 VDD.t345 9.52217
R1372 VDD.n470 VDD.t321 9.52217
R1373 VDD.n470 VDD.t357 9.52217
R1374 VDD.n469 VDD.t146 9.52217
R1375 VDD.n469 VDD.t404 9.52217
R1376 VDD.n74 VDD.t291 9.52217
R1377 VDD.n74 VDD.t349 9.52217
R1378 VDD.n70 VDD.t297 9.52217
R1379 VDD.n70 VDD.t261 9.52217
R1380 VDD.n66 VDD.t226 9.52217
R1381 VDD.n66 VDD.t136 9.52217
R1382 VDD.n62 VDD.t343 9.52217
R1383 VDD.n62 VDD.t398 9.52217
R1384 VDD.n58 VDD.t459 9.52217
R1385 VDD.n58 VDD.t275 9.52217
R1386 VDD.n54 VDD.t445 9.52217
R1387 VDD.n54 VDD.t138 9.52217
R1388 VDD.n50 VDD.t5 9.52217
R1389 VDD.n50 VDD.t142 9.52217
R1390 VDD.n46 VDD.t1 9.52217
R1391 VDD.n46 VDD.t140 9.52217
R1392 VDD.n42 VDD.t426 9.52217
R1393 VDD.n42 VDD.t428 9.52217
R1394 VDD.n38 VDD.t420 9.52217
R1395 VDD.n38 VDD.t422 9.52217
R1396 VDD.n34 VDD.t392 9.52217
R1397 VDD.n34 VDD.t390 9.52217
R1398 VDD.n30 VDD.t329 9.52217
R1399 VDD.n30 VDD.t59 9.52217
R1400 VDD.n26 VDD.t361 9.52217
R1401 VDD.n26 VDD.t367 9.52217
R1402 VDD.n22 VDD.t363 9.52217
R1403 VDD.n22 VDD.t439 9.52217
R1404 VDD.n1 VDD.t223 9.52217
R1405 VDD.n1 VDD.t406 9.52217
R1406 VDD.n4 VDD.t87 9.52217
R1407 VDD.n4 VDD.t503 9.52217
R1408 VDD.n460 VDD.n459 6.60764
R1409 VDD.n450 VDD.n449 6.60764
R1410 VDD.n440 VDD.n439 6.60764
R1411 VDD.n430 VDD.n429 6.60764
R1412 VDD.n420 VDD.n419 6.60764
R1413 VDD.n410 VDD.n409 6.60764
R1414 VDD.n400 VDD.n399 6.60764
R1415 VDD.n391 VDD.n390 6.60764
R1416 VDD.n463 VDD.n459 5.77063
R1417 VDD.n453 VDD.n449 5.77063
R1418 VDD.n443 VDD.n439 5.77063
R1419 VDD.n433 VDD.n429 5.77063
R1420 VDD.n423 VDD.n419 5.77063
R1421 VDD.n413 VDD.n409 5.77063
R1422 VDD.n403 VDD.n399 5.77063
R1423 VDD.n394 VDD.n390 5.77063
R1424 VDD.t446 VDD.n173 5.4667
R1425 VDD.n255 VDD.t160 5.4667
R1426 VDD.t475 VDD.n583 5.4667
R1427 VDD.n605 VDD.t191 5.4667
R1428 VDD.n933 VDD.n72 5.44168
R1429 VDD.n927 VDD.n72 5.44168
R1430 VDD.n947 VDD.n64 5.44168
R1431 VDD.n941 VDD.n64 5.44168
R1432 VDD.n961 VDD.n56 5.44168
R1433 VDD.n955 VDD.n56 5.44168
R1434 VDD.n975 VDD.n48 5.44168
R1435 VDD.n969 VDD.n48 5.44168
R1436 VDD.n989 VDD.n40 5.44168
R1437 VDD.n983 VDD.n40 5.44168
R1438 VDD.n1003 VDD.n32 5.44168
R1439 VDD.n997 VDD.n32 5.44168
R1440 VDD.n1017 VDD.n24 5.44168
R1441 VDD.n1011 VDD.n24 5.44168
R1442 VDD.n15 VDD.n13 5.44168
R1443 VDD.n13 VDD.n12 5.44168
R1444 VDD.n915 VDD.n721 5.0005
R1445 VDD.n900 VDD.n729 5.0005
R1446 VDD.n885 VDD.n737 5.0005
R1447 VDD.n870 VDD.n745 5.0005
R1448 VDD.n855 VDD.n753 5.0005
R1449 VDD.n840 VDD.n761 5.0005
R1450 VDD.n825 VDD.n769 5.0005
R1451 VDD.n810 VDD.n777 5.0005
R1452 VDD.n795 VDD.n785 5.0005
R1453 VDD.n554 VDD.n548 5.0005
R1454 VDD.n541 VDD.n535 5.0005
R1455 VDD.n528 VDD.n522 5.0005
R1456 VDD.n515 VDD.n509 5.0005
R1457 VDD.n502 VDD.n496 5.0005
R1458 VDD.n489 VDD.n483 5.0005
R1459 VDD.n479 VDD.n474 5.0005
R1460 VDD.n914 VDD.n912 3.72599
R1461 VDD.n899 VDD.n897 3.72599
R1462 VDD.n884 VDD.n882 3.72599
R1463 VDD.n869 VDD.n867 3.72599
R1464 VDD.n854 VDD.n852 3.72599
R1465 VDD.n839 VDD.n837 3.72599
R1466 VDD.n824 VDD.n822 3.72599
R1467 VDD.n809 VDD.n807 3.72599
R1468 VDD.n794 VDD.n792 3.72599
R1469 VDD.n482 VDD.n481 3.72599
R1470 VDD.n495 VDD.n494 3.72599
R1471 VDD.n508 VDD.n507 3.72599
R1472 VDD.n521 VDD.n520 3.72599
R1473 VDD.n534 VDD.n533 3.72599
R1474 VDD.n547 VDD.n546 3.72599
R1475 VDD.n640 VDD.n639 3.72599
R1476 VDD VDD.n923 2.86795
R1477 VDD.n6 VDD.n5 2.53478
R1478 VDD.n925 VDD.n72 2.35344
R1479 VDD.n939 VDD.n64 2.35344
R1480 VDD.n953 VDD.n56 2.35344
R1481 VDD.n967 VDD.n48 2.35344
R1482 VDD.n981 VDD.n40 2.35344
R1483 VDD.n995 VDD.n32 2.35344
R1484 VDD.n1009 VDD.n24 2.35344
R1485 VDD.n13 VDD.n8 2.35344
R1486 VDD.n261 VDD.n260 2.3255
R1487 VDD.n264 VDD.n263 2.3255
R1488 VDD.n268 VDD.n267 2.3255
R1489 VDD.n271 VDD.n270 2.3255
R1490 VDD.n275 VDD.n274 2.3255
R1491 VDD.n278 VDD.n277 2.3255
R1492 VDD.n282 VDD.n281 2.3255
R1493 VDD.n285 VDD.n284 2.3255
R1494 VDD.n289 VDD.n288 2.3255
R1495 VDD.n292 VDD.n291 2.3255
R1496 VDD.n296 VDD.n295 2.3255
R1497 VDD.n299 VDD.n298 2.3255
R1498 VDD.n303 VDD.n302 2.3255
R1499 VDD.n306 VDD.n305 2.3255
R1500 VDD.n310 VDD.n309 2.3255
R1501 VDD.n313 VDD.n312 2.3255
R1502 VDD.n317 VDD.n316 2.3255
R1503 VDD.n320 VDD.n319 2.3255
R1504 VDD.n324 VDD.n323 2.3255
R1505 VDD.n327 VDD.n326 2.3255
R1506 VDD.n331 VDD.n330 2.3255
R1507 VDD.n334 VDD.n333 2.3255
R1508 VDD.n338 VDD.n337 2.3255
R1509 VDD.n341 VDD.n340 2.3255
R1510 VDD.n345 VDD.n344 2.3255
R1511 VDD.n348 VDD.n347 2.3255
R1512 VDD.n352 VDD.n351 2.3255
R1513 VDD.n355 VDD.n354 2.3255
R1514 VDD.n611 VDD.n610 2.3255
R1515 VDD.n614 VDD.n613 2.3255
R1516 VDD.n618 VDD.n617 2.3255
R1517 VDD.n621 VDD.n620 2.3255
R1518 VDD.n625 VDD.n624 2.3255
R1519 VDD.n628 VDD.n627 2.3255
R1520 VDD.n632 VDD.n631 2.3255
R1521 VDD.n635 VDD.n634 2.3255
R1522 VDD.n931 VDD.n924 2.29581
R1523 VDD.n73 VDD.n71 2.29581
R1524 VDD.n937 VDD.n69 2.29581
R1525 VDD.n945 VDD.n938 2.29581
R1526 VDD.n65 VDD.n63 2.29581
R1527 VDD.n951 VDD.n61 2.29581
R1528 VDD.n959 VDD.n952 2.29581
R1529 VDD.n57 VDD.n55 2.29581
R1530 VDD.n965 VDD.n53 2.29581
R1531 VDD.n973 VDD.n966 2.29581
R1532 VDD.n49 VDD.n47 2.29581
R1533 VDD.n979 VDD.n45 2.29581
R1534 VDD.n987 VDD.n980 2.29581
R1535 VDD.n41 VDD.n39 2.29581
R1536 VDD.n993 VDD.n37 2.29581
R1537 VDD.n1001 VDD.n994 2.29581
R1538 VDD.n33 VDD.n31 2.29581
R1539 VDD.n1007 VDD.n29 2.29581
R1540 VDD.n1015 VDD.n1008 2.29581
R1541 VDD.n25 VDD.n23 2.29581
R1542 VDD.n1021 VDD.n21 2.29581
R1543 VDD.n20 VDD.n0 2.29581
R1544 VDD.n17 VDD.n2 2.29581
R1545 VDD.n789 VDD.n788 2.1858
R1546 VDD.n83 VDD.n80 2.04321
R1547 VDD.n90 VDD.n87 2.04321
R1548 VDD.n342 VDD.n91 2.04321
R1549 VDD.n97 VDD.n94 2.04321
R1550 VDD.n335 VDD.n98 2.04321
R1551 VDD.n104 VDD.n101 2.04321
R1552 VDD.n328 VDD.n105 2.04321
R1553 VDD.n111 VDD.n108 2.04321
R1554 VDD.n321 VDD.n112 2.04321
R1555 VDD.n118 VDD.n115 2.04321
R1556 VDD.n314 VDD.n119 2.04321
R1557 VDD.n125 VDD.n122 2.04321
R1558 VDD.n307 VDD.n126 2.04321
R1559 VDD.n132 VDD.n129 2.04321
R1560 VDD.n300 VDD.n133 2.04321
R1561 VDD.n139 VDD.n136 2.04321
R1562 VDD.n293 VDD.n140 2.04321
R1563 VDD.n146 VDD.n143 2.04321
R1564 VDD.n286 VDD.n147 2.04321
R1565 VDD.n153 VDD.n150 2.04321
R1566 VDD.n279 VDD.n154 2.04321
R1567 VDD.n160 VDD.n157 2.04321
R1568 VDD.n272 VDD.n161 2.04321
R1569 VDD.n167 VDD.n164 2.04321
R1570 VDD.n265 VDD.n168 2.04321
R1571 VDD.n257 VDD.n171 2.04321
R1572 VDD.n258 VDD.n256 2.04321
R1573 VDD.n349 VDD.n84 2.04321
R1574 VDD.n356 VDD.n77 2.04321
R1575 VDD.n563 VDD.n560 2.04321
R1576 VDD.n570 VDD.n567 2.04321
R1577 VDD.n622 VDD.n571 2.04321
R1578 VDD.n577 VDD.n574 2.04321
R1579 VDD.n615 VDD.n578 2.04321
R1580 VDD.n607 VDD.n581 2.04321
R1581 VDD.n608 VDD.n606 2.04321
R1582 VDD.n629 VDD.n564 2.04321
R1583 VDD.n636 VDD.n557 2.04321
R1584 VDD.n929 VDD.n927 1.97967
R1585 VDD.n943 VDD.n941 1.97967
R1586 VDD.n957 VDD.n955 1.97967
R1587 VDD.n971 VDD.n969 1.97967
R1588 VDD.n985 VDD.n983 1.97967
R1589 VDD.n999 VDD.n997 1.97967
R1590 VDD.n1013 VDD.n1011 1.97967
R1591 VDD.n12 VDD.n11 1.97967
R1592 VDD.n920 VDD.n715 1.9397
R1593 VDD.n909 VDD.n908 1.9397
R1594 VDD.n905 VDD.n723 1.9397
R1595 VDD.n894 VDD.n893 1.9397
R1596 VDD.n890 VDD.n731 1.9397
R1597 VDD.n879 VDD.n878 1.9397
R1598 VDD.n875 VDD.n739 1.9397
R1599 VDD.n864 VDD.n863 1.9397
R1600 VDD.n860 VDD.n747 1.9397
R1601 VDD.n849 VDD.n848 1.9397
R1602 VDD.n845 VDD.n755 1.9397
R1603 VDD.n834 VDD.n833 1.9397
R1604 VDD.n830 VDD.n763 1.9397
R1605 VDD.n819 VDD.n818 1.9397
R1606 VDD.n815 VDD.n771 1.9397
R1607 VDD.n804 VDD.n803 1.9397
R1608 VDD.n800 VDD.n779 1.9397
R1609 VDD.n643 VDD.n637 1.9397
R1610 VDD.n649 VDD.n648 1.9397
R1611 VDD.n654 VDD.n544 1.9397
R1612 VDD.n660 VDD.n659 1.9397
R1613 VDD.n665 VDD.n531 1.9397
R1614 VDD.n671 VDD.n670 1.9397
R1615 VDD.n676 VDD.n518 1.9397
R1616 VDD.n682 VDD.n681 1.9397
R1617 VDD.n687 VDD.n505 1.9397
R1618 VDD.n693 VDD.n692 1.9397
R1619 VDD.n698 VDD.n492 1.9397
R1620 VDD.n704 VDD.n703 1.9397
R1621 VDD.n709 VDD.n477 1.9397
R1622 VDD.n714 VDD.n468 1.9397
R1623 VDD.n467 VDD.n357 1.91627
R1624 VDD.n457 VDD.n361 1.91627
R1625 VDD.n447 VDD.n365 1.91627
R1626 VDD.n437 VDD.n369 1.91627
R1627 VDD.n427 VDD.n373 1.91627
R1628 VDD.n417 VDD.n377 1.91627
R1629 VDD.n407 VDD.n381 1.91627
R1630 VDD.n397 VDD.n385 1.91627
R1631 VDD.n803 VDD.n800 1.52654
R1632 VDD.n818 VDD.n815 1.52654
R1633 VDD.n833 VDD.n830 1.52654
R1634 VDD.n848 VDD.n845 1.52654
R1635 VDD.n863 VDD.n860 1.52654
R1636 VDD.n878 VDD.n875 1.52654
R1637 VDD.n893 VDD.n890 1.52654
R1638 VDD.n908 VDD.n905 1.52654
R1639 VDD.n922 VDD 1.42472
R1640 VDD.n405 VDD 1.04243
R1641 VDD.n415 VDD 1.04243
R1642 VDD.n425 VDD 1.04243
R1643 VDD.n435 VDD 1.04243
R1644 VDD.n445 VDD 1.04243
R1645 VDD.n455 VDD 1.04243
R1646 VDD.n465 VDD 1.04243
R1647 VDD.n359 VDD.n358 0.957022
R1648 VDD.n363 VDD.n362 0.957022
R1649 VDD.n367 VDD.n366 0.957022
R1650 VDD.n371 VDD.n370 0.957022
R1651 VDD.n375 VDD.n374 0.957022
R1652 VDD.n379 VDD.n378 0.957022
R1653 VDD.n383 VDD.n382 0.957022
R1654 VDD.n387 VDD.n386 0.957022
R1655 VDD.n923 VDD.n356 0.948417
R1656 VDD.n921 VDD.n920 0.727062
R1657 VDD.n464 VDD.n463 0.713588
R1658 VDD.n454 VDD.n453 0.713588
R1659 VDD.n444 VDD.n443 0.713588
R1660 VDD.n434 VDD.n433 0.713588
R1661 VDD.n424 VDD.n423 0.713588
R1662 VDD.n414 VDD.n413 0.713588
R1663 VDD.n404 VDD.n403 0.713588
R1664 VDD.n395 VDD.n394 0.713588
R1665 VDD VDD.n1021 0.669618
R1666 VDD VDD.n1007 0.669618
R1667 VDD VDD.n993 0.669618
R1668 VDD VDD.n979 0.669618
R1669 VDD VDD.n965 0.669618
R1670 VDD VDD.n951 0.669618
R1671 VDD VDD.n937 0.669618
R1672 VDD.n396 VDD.n395 0.647749
R1673 VDD.n711 VDD.n710 0.6205
R1674 VDD.n700 VDD.n699 0.6205
R1675 VDD.n689 VDD.n688 0.6205
R1676 VDD.n678 VDD.n677 0.6205
R1677 VDD.n667 VDD.n666 0.6205
R1678 VDD.n656 VDD.n655 0.6205
R1679 VDD.n645 VDD.n644 0.6205
R1680 VDD.n797 VDD.n796 0.6205
R1681 VDD.n812 VDD.n811 0.6205
R1682 VDD.n827 VDD.n826 0.6205
R1683 VDD.n842 VDD.n841 0.6205
R1684 VDD.n857 VDD.n856 0.6205
R1685 VDD.n872 VDD.n871 0.6205
R1686 VDD.n887 VDD.n886 0.6205
R1687 VDD.n902 VDD.n901 0.6205
R1688 VDD.n917 VDD.n916 0.6205
R1689 VDD.n16 VDD.n15 0.58175
R1690 VDD.n1018 VDD.n1017 0.58175
R1691 VDD.n1004 VDD.n1003 0.58175
R1692 VDD.n990 VDD.n989 0.58175
R1693 VDD.n976 VDD.n975 0.58175
R1694 VDD.n962 VDD.n961 0.58175
R1695 VDD.n948 VDD.n947 0.58175
R1696 VDD.n934 VDD.n933 0.58175
R1697 VDD.n916 VDD.n720 0.533833
R1698 VDD.n901 VDD.n728 0.533833
R1699 VDD.n886 VDD.n736 0.533833
R1700 VDD.n871 VDD.n744 0.533833
R1701 VDD.n856 VDD.n752 0.533833
R1702 VDD.n841 VDD.n760 0.533833
R1703 VDD.n826 VDD.n768 0.533833
R1704 VDD.n811 VDD.n776 0.533833
R1705 VDD.n796 VDD.n784 0.533833
R1706 VDD.n644 VDD.n549 0.533833
R1707 VDD.n655 VDD.n536 0.533833
R1708 VDD.n666 VDD.n523 0.533833
R1709 VDD.n677 VDD.n510 0.533833
R1710 VDD.n688 VDD.n497 0.533833
R1711 VDD.n699 VDD.n484 0.533833
R1712 VDD.n710 VDD.n473 0.533833
R1713 VDD.n921 VDD.n714 0.495292
R1714 VDD.n360 VDD.n359 0.478761
R1715 VDD.n364 VDD.n363 0.478761
R1716 VDD.n368 VDD.n367 0.478761
R1717 VDD.n372 VDD.n371 0.478761
R1718 VDD.n376 VDD.n375 0.478761
R1719 VDD.n380 VDD.n379 0.478761
R1720 VDD.n384 VDD.n383 0.478761
R1721 VDD.n388 VDD.n387 0.478761
R1722 VDD VDD.n636 0.438
R1723 VDD VDD.n397 0.394487
R1724 VDD VDD.n407 0.394487
R1725 VDD VDD.n417 0.394487
R1726 VDD VDD.n427 0.394487
R1727 VDD VDD.n437 0.394487
R1728 VDD VDD.n447 0.394487
R1729 VDD VDD.n457 0.394487
R1730 VDD VDD.n467 0.394487
R1731 VDD.n405 VDD.n404 0.358192
R1732 VDD.n415 VDD.n414 0.358192
R1733 VDD.n425 VDD.n424 0.358192
R1734 VDD.n435 VDD.n434 0.358192
R1735 VDD.n445 VDD.n444 0.358192
R1736 VDD.n455 VDD.n454 0.358192
R1737 VDD.n465 VDD.n464 0.358192
R1738 VDD.n922 VDD 0.350184
R1739 VDD.n466 VDD.n360 0.337457
R1740 VDD.n456 VDD.n364 0.337457
R1741 VDD.n446 VDD.n368 0.337457
R1742 VDD.n436 VDD.n372 0.337457
R1743 VDD.n426 VDD.n376 0.337457
R1744 VDD.n416 VDD.n380 0.337457
R1745 VDD.n406 VDD.n384 0.337457
R1746 VDD.n396 VDD.n388 0.337457
R1747 VDD.n5 VDD.n3 0.324029
R1748 VDD.n19 VDD.n18 0.324029
R1749 VDD.n1020 VDD.n1019 0.324029
R1750 VDD.n28 VDD.n27 0.324029
R1751 VDD.n1006 VDD.n1005 0.324029
R1752 VDD.n36 VDD.n35 0.324029
R1753 VDD.n992 VDD.n991 0.324029
R1754 VDD.n44 VDD.n43 0.324029
R1755 VDD.n978 VDD.n977 0.324029
R1756 VDD.n52 VDD.n51 0.324029
R1757 VDD.n964 VDD.n963 0.324029
R1758 VDD.n60 VDD.n59 0.324029
R1759 VDD.n950 VDD.n949 0.324029
R1760 VDD.n68 VDD.n67 0.324029
R1761 VDD.n936 VDD.n935 0.324029
R1762 VDD.n76 VDD.n75 0.324029
R1763 VDD.n406 VDD.n405 0.290057
R1764 VDD.n416 VDD.n415 0.290057
R1765 VDD.n426 VDD.n425 0.290057
R1766 VDD.n436 VDD.n435 0.290057
R1767 VDD.n446 VDD.n445 0.290057
R1768 VDD.n456 VDD.n455 0.290057
R1769 VDD.n466 VDD.n465 0.290057
R1770 VDD.n923 VDD.n922 0.274719
R1771 VDD.n712 VDD.n711 0.253104
R1772 VDD.n701 VDD.n700 0.253104
R1773 VDD.n690 VDD.n689 0.253104
R1774 VDD.n679 VDD.n678 0.253104
R1775 VDD.n668 VDD.n667 0.253104
R1776 VDD.n657 VDD.n656 0.253104
R1777 VDD.n646 VDD.n645 0.253104
R1778 VDD.n797 VDD.n783 0.253104
R1779 VDD.n812 VDD.n775 0.253104
R1780 VDD.n827 VDD.n767 0.253104
R1781 VDD.n842 VDD.n759 0.253104
R1782 VDD.n857 VDD.n751 0.253104
R1783 VDD.n872 VDD.n743 0.253104
R1784 VDD.n887 VDD.n735 0.253104
R1785 VDD.n902 VDD.n727 0.253104
R1786 VDD.n917 VDD.n719 0.253104
R1787 VDD.n933 VDD.n932 0.25148
R1788 VDD.n947 VDD.n946 0.25148
R1789 VDD.n961 VDD.n960 0.25148
R1790 VDD.n975 VDD.n974 0.25148
R1791 VDD.n989 VDD.n988 0.25148
R1792 VDD.n1003 VDD.n1002 0.25148
R1793 VDD.n1017 VDD.n1016 0.25148
R1794 VDD.n15 VDD.n14 0.25148
R1795 VDD.n714 VDD.n713 0.246594
R1796 VDD.n477 VDD.n476 0.246594
R1797 VDD.n703 VDD.n702 0.246594
R1798 VDD.n492 VDD.n491 0.246594
R1799 VDD.n692 VDD.n691 0.246594
R1800 VDD.n505 VDD.n504 0.246594
R1801 VDD.n681 VDD.n680 0.246594
R1802 VDD.n518 VDD.n517 0.246594
R1803 VDD.n670 VDD.n669 0.246594
R1804 VDD.n531 VDD.n530 0.246594
R1805 VDD.n659 VDD.n658 0.246594
R1806 VDD.n544 VDD.n543 0.246594
R1807 VDD.n648 VDD.n647 0.246594
R1808 VDD.n637 VDD.n556 0.246594
R1809 VDD.n800 VDD.n799 0.246594
R1810 VDD.n803 VDD.n802 0.246594
R1811 VDD.n815 VDD.n814 0.246594
R1812 VDD.n818 VDD.n817 0.246594
R1813 VDD.n830 VDD.n829 0.246594
R1814 VDD.n833 VDD.n832 0.246594
R1815 VDD.n845 VDD.n844 0.246594
R1816 VDD.n848 VDD.n847 0.246594
R1817 VDD.n860 VDD.n859 0.246594
R1818 VDD.n863 VDD.n862 0.246594
R1819 VDD.n875 VDD.n874 0.246594
R1820 VDD.n878 VDD.n877 0.246594
R1821 VDD.n890 VDD.n889 0.246594
R1822 VDD.n893 VDD.n892 0.246594
R1823 VDD.n905 VDD.n904 0.246594
R1824 VDD.n908 VDD.n907 0.246594
R1825 VDD.n920 VDD.n919 0.246594
R1826 VDD.n711 VDD.n472 0.242688
R1827 VDD.n700 VDD.n488 0.242688
R1828 VDD.n689 VDD.n501 0.242688
R1829 VDD.n678 VDD.n514 0.242688
R1830 VDD.n667 VDD.n527 0.242688
R1831 VDD.n656 VDD.n540 0.242688
R1832 VDD.n645 VDD.n553 0.242688
R1833 VDD.n798 VDD.n797 0.242688
R1834 VDD.n813 VDD.n812 0.242688
R1835 VDD.n828 VDD.n827 0.242688
R1836 VDD.n843 VDD.n842 0.242688
R1837 VDD.n858 VDD.n857 0.242688
R1838 VDD.n873 VDD.n872 0.242688
R1839 VDD.n888 VDD.n887 0.242688
R1840 VDD.n903 VDD.n902 0.242688
R1841 VDD.n918 VDD.n917 0.242688
R1842 VDD.n1021 VDD.n1020 0.239471
R1843 VDD.n1007 VDD.n1006 0.239471
R1844 VDD.n993 VDD.n992 0.239471
R1845 VDD.n979 VDD.n978 0.239471
R1846 VDD.n965 VDD.n964 0.239471
R1847 VDD.n951 VDD.n950 0.239471
R1848 VDD.n937 VDD.n936 0.239471
R1849 VDD.n20 VDD.n19 0.232118
R1850 VDD.n1008 VDD.n28 0.232118
R1851 VDD.n994 VDD.n36 0.232118
R1852 VDD.n980 VDD.n44 0.232118
R1853 VDD.n966 VDD.n52 0.232118
R1854 VDD.n952 VDD.n60 0.232118
R1855 VDD.n938 VDD.n68 0.232118
R1856 VDD.n924 VDD.n76 0.232118
R1857 VDD.n713 VDD.n712 0.229667
R1858 VDD.n476 VDD.n472 0.229667
R1859 VDD.n702 VDD.n701 0.229667
R1860 VDD.n491 VDD.n488 0.229667
R1861 VDD.n691 VDD.n690 0.229667
R1862 VDD.n504 VDD.n501 0.229667
R1863 VDD.n680 VDD.n679 0.229667
R1864 VDD.n517 VDD.n514 0.229667
R1865 VDD.n669 VDD.n668 0.229667
R1866 VDD.n530 VDD.n527 0.229667
R1867 VDD.n658 VDD.n657 0.229667
R1868 VDD.n543 VDD.n540 0.229667
R1869 VDD.n647 VDD.n646 0.229667
R1870 VDD.n556 VDD.n553 0.229667
R1871 VDD.n788 VDD.n783 0.229667
R1872 VDD.n799 VDD.n798 0.229667
R1873 VDD.n802 VDD.n775 0.229667
R1874 VDD.n814 VDD.n813 0.229667
R1875 VDD.n817 VDD.n767 0.229667
R1876 VDD.n829 VDD.n828 0.229667
R1877 VDD.n832 VDD.n759 0.229667
R1878 VDD.n844 VDD.n843 0.229667
R1879 VDD.n847 VDD.n751 0.229667
R1880 VDD.n859 VDD.n858 0.229667
R1881 VDD.n862 VDD.n743 0.229667
R1882 VDD.n874 VDD.n873 0.229667
R1883 VDD.n877 VDD.n735 0.229667
R1884 VDD.n889 VDD.n888 0.229667
R1885 VDD.n892 VDD.n727 0.229667
R1886 VDD.n904 VDD.n903 0.229667
R1887 VDD.n907 VDD.n719 0.229667
R1888 VDD.n919 VDD.n918 0.229667
R1889 VDD.n703 VDD.n477 0.221854
R1890 VDD.n692 VDD.n492 0.221854
R1891 VDD.n681 VDD.n505 0.221854
R1892 VDD.n670 VDD.n518 0.221854
R1893 VDD.n659 VDD.n531 0.221854
R1894 VDD.n648 VDD.n544 0.221854
R1895 VDD.n356 VDD.n355 0.189302
R1896 VDD.n351 VDD.n83 0.189302
R1897 VDD.n349 VDD.n348 0.189302
R1898 VDD.n344 VDD.n90 0.189302
R1899 VDD.n342 VDD.n341 0.189302
R1900 VDD.n337 VDD.n97 0.189302
R1901 VDD.n335 VDD.n334 0.189302
R1902 VDD.n330 VDD.n104 0.189302
R1903 VDD.n328 VDD.n327 0.189302
R1904 VDD.n323 VDD.n111 0.189302
R1905 VDD.n321 VDD.n320 0.189302
R1906 VDD.n316 VDD.n118 0.189302
R1907 VDD.n314 VDD.n313 0.189302
R1908 VDD.n309 VDD.n125 0.189302
R1909 VDD.n307 VDD.n306 0.189302
R1910 VDD.n302 VDD.n132 0.189302
R1911 VDD.n300 VDD.n299 0.189302
R1912 VDD.n295 VDD.n139 0.189302
R1913 VDD.n293 VDD.n292 0.189302
R1914 VDD.n288 VDD.n146 0.189302
R1915 VDD.n286 VDD.n285 0.189302
R1916 VDD.n281 VDD.n153 0.189302
R1917 VDD.n279 VDD.n278 0.189302
R1918 VDD.n274 VDD.n160 0.189302
R1919 VDD.n272 VDD.n271 0.189302
R1920 VDD.n267 VDD.n167 0.189302
R1921 VDD.n265 VDD.n264 0.189302
R1922 VDD.n260 VDD.n257 0.189302
R1923 VDD.n636 VDD.n635 0.189302
R1924 VDD.n631 VDD.n563 0.189302
R1925 VDD.n629 VDD.n628 0.189302
R1926 VDD.n624 VDD.n570 0.189302
R1927 VDD.n622 VDD.n621 0.189302
R1928 VDD.n617 VDD.n577 0.189302
R1929 VDD.n615 VDD.n614 0.189302
R1930 VDD.n610 VDD.n607 0.189302
R1931 VDD.n637 VDD 0.151542
R1932 VDD.n83 VDD.n78 0.13201
R1933 VDD.n350 VDD.n349 0.13201
R1934 VDD.n90 VDD.n85 0.13201
R1935 VDD.n343 VDD.n342 0.13201
R1936 VDD.n97 VDD.n92 0.13201
R1937 VDD.n336 VDD.n335 0.13201
R1938 VDD.n104 VDD.n99 0.13201
R1939 VDD.n329 VDD.n328 0.13201
R1940 VDD.n111 VDD.n106 0.13201
R1941 VDD.n322 VDD.n321 0.13201
R1942 VDD.n118 VDD.n113 0.13201
R1943 VDD.n315 VDD.n314 0.13201
R1944 VDD.n125 VDD.n120 0.13201
R1945 VDD.n308 VDD.n307 0.13201
R1946 VDD.n132 VDD.n127 0.13201
R1947 VDD.n301 VDD.n300 0.13201
R1948 VDD.n139 VDD.n134 0.13201
R1949 VDD.n294 VDD.n293 0.13201
R1950 VDD.n146 VDD.n141 0.13201
R1951 VDD.n287 VDD.n286 0.13201
R1952 VDD.n153 VDD.n148 0.13201
R1953 VDD.n280 VDD.n279 0.13201
R1954 VDD.n160 VDD.n155 0.13201
R1955 VDD.n273 VDD.n272 0.13201
R1956 VDD.n167 VDD.n162 0.13201
R1957 VDD.n266 VDD.n265 0.13201
R1958 VDD.n257 VDD.n169 0.13201
R1959 VDD.n259 VDD.n258 0.13201
R1960 VDD.n563 VDD.n558 0.13201
R1961 VDD.n630 VDD.n629 0.13201
R1962 VDD.n570 VDD.n565 0.13201
R1963 VDD.n623 VDD.n622 0.13201
R1964 VDD.n577 VDD.n572 0.13201
R1965 VDD.n616 VDD.n615 0.13201
R1966 VDD.n607 VDD.n579 0.13201
R1967 VDD.n609 VDD.n608 0.13201
R1968 VDD.n18 VDD.n17 0.124275
R1969 VDD.n27 VDD.n23 0.124275
R1970 VDD.n35 VDD.n31 0.124275
R1971 VDD.n43 VDD.n39 0.124275
R1972 VDD.n51 VDD.n47 0.124275
R1973 VDD.n59 VDD.n55 0.124275
R1974 VDD.n67 VDD.n63 0.124275
R1975 VDD.n75 VDD.n71 0.124275
R1976 VDD.n16 VDD.n3 0.121824
R1977 VDD.n1019 VDD.n1018 0.121824
R1978 VDD.n1005 VDD.n1004 0.121824
R1979 VDD.n991 VDD.n990 0.121824
R1980 VDD.n977 VDD.n976 0.121824
R1981 VDD.n963 VDD.n962 0.121824
R1982 VDD.n949 VDD.n948 0.121824
R1983 VDD.n935 VDD.n934 0.121824
R1984 VDD VDD.n20 0.113245
R1985 VDD.n1008 VDD 0.113245
R1986 VDD.n994 VDD 0.113245
R1987 VDD.n980 VDD 0.113245
R1988 VDD.n966 VDD 0.113245
R1989 VDD.n952 VDD 0.113245
R1990 VDD.n938 VDD 0.113245
R1991 VDD.n924 VDD 0.113245
R1992 VDD.n397 VDD.n396 0.0804051
R1993 VDD.n407 VDD.n406 0.0804051
R1994 VDD.n417 VDD.n416 0.0804051
R1995 VDD.n427 VDD.n426 0.0804051
R1996 VDD.n437 VDD.n436 0.0804051
R1997 VDD.n447 VDD.n446 0.0804051
R1998 VDD.n457 VDD.n456 0.0804051
R1999 VDD.n467 VDD.n466 0.0804051
R2000 VDD.n258 VDD 0.0708125
R2001 VDD.n608 VDD 0.0708125
R2002 VDD.n355 VDD.n78 0.0577917
R2003 VDD.n351 VDD.n350 0.0577917
R2004 VDD.n348 VDD.n85 0.0577917
R2005 VDD.n344 VDD.n343 0.0577917
R2006 VDD.n341 VDD.n92 0.0577917
R2007 VDD.n337 VDD.n336 0.0577917
R2008 VDD.n334 VDD.n99 0.0577917
R2009 VDD.n330 VDD.n329 0.0577917
R2010 VDD.n327 VDD.n106 0.0577917
R2011 VDD.n323 VDD.n322 0.0577917
R2012 VDD.n320 VDD.n113 0.0577917
R2013 VDD.n316 VDD.n315 0.0577917
R2014 VDD.n313 VDD.n120 0.0577917
R2015 VDD.n309 VDD.n308 0.0577917
R2016 VDD.n306 VDD.n127 0.0577917
R2017 VDD.n302 VDD.n301 0.0577917
R2018 VDD.n299 VDD.n134 0.0577917
R2019 VDD.n295 VDD.n294 0.0577917
R2020 VDD.n292 VDD.n141 0.0577917
R2021 VDD.n288 VDD.n287 0.0577917
R2022 VDD.n285 VDD.n148 0.0577917
R2023 VDD.n281 VDD.n280 0.0577917
R2024 VDD.n278 VDD.n155 0.0577917
R2025 VDD.n274 VDD.n273 0.0577917
R2026 VDD.n271 VDD.n162 0.0577917
R2027 VDD.n267 VDD.n266 0.0577917
R2028 VDD.n264 VDD.n169 0.0577917
R2029 VDD.n260 VDD.n259 0.0577917
R2030 VDD.n635 VDD.n558 0.0577917
R2031 VDD.n631 VDD.n630 0.0577917
R2032 VDD.n628 VDD.n565 0.0577917
R2033 VDD.n624 VDD.n623 0.0577917
R2034 VDD.n621 VDD.n572 0.0577917
R2035 VDD.n617 VDD.n616 0.0577917
R2036 VDD.n614 VDD.n579 0.0577917
R2037 VDD.n610 VDD.n609 0.0577917
R2038 VDD VDD.n921 0.013
R2039 VDD.n17 VDD.n16 0.00295098
R2040 VDD.n1018 VDD.n23 0.00295098
R2041 VDD.n1004 VDD.n31 0.00295098
R2042 VDD.n990 VDD.n39 0.00295098
R2043 VDD.n976 VDD.n47 0.00295098
R2044 VDD.n962 VDD.n55 0.00295098
R2045 VDD.n948 VDD.n63 0.00295098
R2046 VDD.n934 VDD.n71 0.00295098
R2047 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 879.481
R2048 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 742.783
R2049 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 665.16
R2050 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 623.388
R2051 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 523.774
R2052 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 431.807
R2053 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 427.875
R2054 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 357.26
R2055 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 208.537
R2056 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 168.077
R2057 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R2058 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R2059 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R2060 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 11.1806
R2061 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R2062 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R2063 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R2064 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R2065 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R2066 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 890.727
R2067 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 742.783
R2068 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 665.16
R2069 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 623.388
R2070 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 523.774
R2071 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 431.807
R2072 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 427.875
R2073 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 364.733
R2074 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 208.5
R2075 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 168.007
R2076 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R2077 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 31.2728
R2078 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R2079 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R2080 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R2081 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R2082 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 8.00471
R2083 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R2084 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R2085 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R2086 term_7.n1 term_7.t5 734.539
R2087 term_7.n1 term_7.t4 233.26
R2088 term_7.n2 term_7.n1 162.399
R2089 term_7.n2 term_7.n0 75.5108
R2090 term_7.n4 term_7.n3 66.3172
R2091 term_7.n3 term_7.t3 17.4005
R2092 term_7.n3 term_7.t1 17.4005
R2093 term_7.n0 term_7.t0 9.52217
R2094 term_7.n0 term_7.t2 9.52217
R2095 term_7 term_7.n4 5.08746
R2096 term_7.n4 term_7.n2 0.3755
R2097 VSS.n554 VSS.n114 133481
R2098 VSS.t537 VSS.n554 58429.2
R2099 VSS.n799 VSS.n752 31435.8
R2100 VSS.n752 VSS.n751 29666.5
R2101 VSS.n832 VSS.n752 22512.6
R2102 VSS.n554 VSS.t424 22478
R2103 VSS.n113 VSS.n56 18773.3
R2104 VSS.n946 VSS.n56 18773.3
R2105 VSS.n946 VSS.n34 18773.3
R2106 VSS.n1024 VSS.n34 18773.3
R2107 VSS.n1024 VSS.n12 18773.3
R2108 VSS.n751 VSS.n12 18773.3
R2109 VSS.n114 VSS.n113 18773.3
R2110 VSS.t18 VSS.t16 7780.49
R2111 VSS.n1158 VSS.n636 5774.44
R2112 VSS.n1147 VSS.n651 5774.44
R2113 VSS.n1136 VSS.n666 5774.44
R2114 VSS.n1125 VSS.n681 5774.44
R2115 VSS.n1114 VSS.n696 5774.44
R2116 VSS.n1103 VSS.n711 5774.44
R2117 VSS.n1092 VSS.n1091 5774.44
R2118 VSS.n626 VSS.n114 5547.41
R2119 VSS.n633 VSS.n113 5137.73
R2120 VSS.n1198 VSS.n56 5137.73
R2121 VSS.n947 VSS.n946 5137.73
R2122 VSS.n1216 VSS.n34 5137.73
R2123 VSS.n1025 VSS.n1024 5137.73
R2124 VSS.n1234 VSS.n12 5137.73
R2125 VSS.n751 VSS.n750 5137.73
R2126 VSS.n1169 VSS.n1168 4338.44
R2127 VSS.n912 VSS.n904 4042.48
R2128 VSS.n956 VSS.n938 4042.48
R2129 VSS.n990 VSS.n982 4042.48
R2130 VSS.n1034 VSS.n1016 4042.48
R2131 VSS.n1068 VSS.n1060 4042.48
R2132 VSS.n857 VSS.n855 4042.48
R2133 VSS.n90 VSS.n89 4042.48
R2134 VSS.n835 VSS.n744 4042.48
R2135 VSS.n1199 VSS.n55 3781.58
R2136 VSS.n949 VSS.n948 3781.58
R2137 VSS.n1217 VSS.n33 3781.58
R2138 VSS.n1027 VSS.n1026 3781.58
R2139 VSS.n1235 VSS.n11 3781.58
R2140 VSS.n1090 VSS.n728 3781.58
R2141 VSS.n635 VSS.n634 3781.58
R2142 VSS.n827 VSS.n752 3648.24
R2143 VSS.n912 VSS.n911 3140.17
R2144 VSS.n956 VSS.n955 3140.17
R2145 VSS.n990 VSS.n989 3140.17
R2146 VSS.n1034 VSS.n1033 3140.17
R2147 VSS.n1068 VSS.n1067 3140.17
R2148 VSS.n864 VSS.n857 3140.17
R2149 VSS.n104 VSS.n90 3140.17
R2150 VSS.n835 VSS.n834 3140.17
R2151 VSS.n921 VSS.n897 3120.05
R2152 VSS.n965 VSS.n931 3120.05
R2153 VSS.n999 VSS.n975 3120.05
R2154 VSS.n1043 VSS.n1009 3120.05
R2155 VSS.n1077 VSS.n1053 3120.05
R2156 VSS.n874 VSS.n730 3120.05
R2157 VSS.n1178 VSS.n82 3120.05
R2158 VSS.n843 VSS.n737 3120.05
R2159 VSS.n1198 VSS.n1197 3093.4
R2160 VSS.n947 VSS.n945 3093.4
R2161 VSS.n1216 VSS.n1215 3093.4
R2162 VSS.n1025 VSS.n1023 3093.4
R2163 VSS.n1234 VSS.n1233 3093.4
R2164 VSS.n750 VSS.n749 3093.4
R2165 VSS.n633 VSS.n632 3093.4
R2166 VSS.n802 VSS.n801 3092.2
R2167 VSS.n627 VSS.n91 2755.48
R2168 VSS.n921 VSS.n896 2350.81
R2169 VSS.n965 VSS.n930 2350.81
R2170 VSS.n999 VSS.n974 2350.81
R2171 VSS.n1043 VSS.n1008 2350.81
R2172 VSS.n1077 VSS.n1052 2350.81
R2173 VSS.n1088 VSS.n730 2350.81
R2174 VSS.n1178 VSS.n81 2350.81
R2175 VSS.n843 VSS.n736 2350.81
R2176 VSS.n567 VSS.n566 2227.12
R2177 VSS.n1170 VSS.n1169 2195.13
R2178 VSS.n807 VSS.n786 2099.08
R2179 VSS.n1097 VSS.n725 2099.08
R2180 VSS.n1108 VSS.n710 2099.08
R2181 VSS.n1119 VSS.n695 2099.08
R2182 VSS.n1130 VSS.n680 2099.08
R2183 VSS.n1141 VSS.n665 2099.08
R2184 VSS.n1152 VSS.n650 2099.08
R2185 VSS.n1163 VSS.n102 2099.08
R2186 VSS.n797 VSS.n796 2093.29
R2187 VSS.n1101 VSS.n712 2093.29
R2188 VSS.n1112 VSS.n697 2093.29
R2189 VSS.n1123 VSS.n682 2093.29
R2190 VSS.n1134 VSS.n667 2093.29
R2191 VSS.n1145 VSS.n652 2093.29
R2192 VSS.n1156 VSS.n637 2093.29
R2193 VSS.n1167 VSS.n93 2093.29
R2194 VSS.n511 VSS.n180 2058.56
R2195 VSS.n585 VSS.n180 2058.56
R2196 VSS.n588 VSS.n173 2058.56
R2197 VSS.n177 VSS.n173 2058.56
R2198 VSS.n175 VSS.n154 2058.56
R2199 VSS.n601 VSS.n154 2058.56
R2200 VSS.n604 VSS.n147 2058.56
R2201 VSS.n151 VSS.n147 2058.56
R2202 VSS.n149 VSS.n128 2058.56
R2203 VSS.n617 VSS.n128 2058.56
R2204 VSS.n624 VSS.n115 2058.56
R2205 VSS.n620 VSS.n115 2058.56
R2206 VSS.n513 VSS.n196 2058.56
R2207 VSS.n514 VSS.n513 2058.56
R2208 VSS.n825 VSS.n753 2058.56
R2209 VSS.n798 VSS.n753 2058.56
R2210 VSS.n748 VSS.n10 2058.56
R2211 VSS.n1237 VSS.n10 2058.56
R2212 VSS.n1022 VSS.n32 2058.56
R2213 VSS.n1219 VSS.n32 2058.56
R2214 VSS.n944 VSS.n54 2058.56
R2215 VSS.n1201 VSS.n54 2058.56
R2216 VSS.n111 VSS.n57 2058.56
R2217 VSS.n1196 VSS.n57 2058.56
R2218 VSS.n941 VSS.n35 2058.56
R2219 VSS.n1214 VSS.n35 2058.56
R2220 VSS.n1019 VSS.n13 2058.56
R2221 VSS.n1232 VSS.n13 2058.56
R2222 VSS.n766 VSS.n763 2058.56
R2223 VSS.n763 VSS.n762 2058.56
R2224 VSS.n630 VSS.n73 2058.56
R2225 VSS.n631 VSS.n630 2058.56
R2226 VSS.n915 VSS.n912 1915.82
R2227 VSS.n959 VSS.n956 1915.82
R2228 VSS.n993 VSS.n990 1915.82
R2229 VSS.n1037 VSS.n1034 1915.82
R2230 VSS.n1071 VSS.n1068 1915.82
R2231 VSS.n871 VSS.n857 1915.82
R2232 VSS.n1172 VSS.n90 1915.82
R2233 VSS.n837 VSS.n835 1915.82
R2234 VSS.n915 VSS.n900 1832.1
R2235 VSS.n959 VSS.n934 1832.1
R2236 VSS.n993 VSS.n978 1832.1
R2237 VSS.n1037 VSS.n1012 1832.1
R2238 VSS.n1071 VSS.n1056 1832.1
R2239 VSS.n871 VSS.n858 1832.1
R2240 VSS.n1172 VSS.n85 1832.1
R2241 VSS.n837 VSS.n740 1832.1
R2242 VSS.n1199 VSS.n1198 1809.14
R2243 VSS.n948 VSS.n947 1809.14
R2244 VSS.n1217 VSS.n1216 1809.14
R2245 VSS.n1026 VSS.n1025 1809.14
R2246 VSS.n1235 VSS.n1234 1809.14
R2247 VSS.n750 VSS.n728 1809.14
R2248 VSS.n634 VSS.n633 1809.14
R2249 VSS.n1200 VSS.n1199 1630.46
R2250 VSS.n948 VSS.n942 1630.46
R2251 VSS.n1218 VSS.n1217 1630.46
R2252 VSS.n1026 VSS.n1020 1630.46
R2253 VSS.n1236 VSS.n1235 1630.46
R2254 VSS.n765 VSS.n728 1630.46
R2255 VSS.n634 VSS.n112 1630.46
R2256 VSS.n908 VSS.n896 1562.99
R2257 VSS.n952 VSS.n930 1562.99
R2258 VSS.n986 VSS.n974 1562.99
R2259 VSS.n1030 VSS.n1008 1562.99
R2260 VSS.n1064 VSS.n1052 1562.99
R2261 VSS.n1088 VSS.n729 1562.99
R2262 VSS.n107 VSS.n81 1562.99
R2263 VSS.n830 VSS.n736 1562.99
R2264 VSS.n628 VSS.n627 1263.93
R2265 VSS.n626 VSS.n625 1228.29
R2266 VSS.n919 VSS.n899 1226.74
R2267 VSS.n963 VSS.n933 1226.74
R2268 VSS.n997 VSS.n977 1226.74
R2269 VSS.n1041 VSS.n1011 1226.74
R2270 VSS.n1075 VSS.n1055 1226.74
R2271 VSS.n867 VSS.n861 1226.74
R2272 VSS.n1176 VSS.n84 1226.74
R2273 VSS.n841 VSS.n739 1226.74
R2274 VSS.n904 VSS.n900 1068.72
R2275 VSS.n938 VSS.n934 1068.72
R2276 VSS.n982 VSS.n978 1068.72
R2277 VSS.n1016 VSS.n1012 1068.72
R2278 VSS.n1060 VSS.n1056 1068.72
R2279 VSS.n858 VSS.n855 1068.72
R2280 VSS.n89 VSS.n85 1068.72
R2281 VSS.n744 VSS.n740 1068.72
R2282 VSS.n535 VSS.n519 1058.19
R2283 VSS.n300 VSS.n299 1058.19
R2284 VSS.n568 VSS.n202 1058.19
R2285 VSS.n804 VSS.n797 1023.31
R2286 VSS.n1094 VSS.n712 1023.31
R2287 VSS.n1105 VSS.n697 1023.31
R2288 VSS.n1116 VSS.n682 1023.31
R2289 VSS.n1127 VSS.n667 1023.31
R2290 VSS.n1138 VSS.n652 1023.31
R2291 VSS.n1149 VSS.n637 1023.31
R2292 VSS.n1160 VSS.n93 1023.31
R2293 VSS.t262 VSS.n1159 994.611
R2294 VSS.t343 VSS.n1148 994.611
R2295 VSS.t419 VSS.n1137 994.611
R2296 VSS.t0 VSS.n1126 994.611
R2297 VSS.t470 VSS.n1115 994.611
R2298 VSS.t112 VSS.n1104 994.611
R2299 VSS.t387 VSS.n1093 994.611
R2300 VSS.t378 VSS.n802 994.611
R2301 VSS.n518 VSS.n517 979.467
R2302 VSS.n1161 VSS.t260 955.091
R2303 VSS.n1168 VSS.t371 955.091
R2304 VSS.n1150 VSS.t305 955.091
R2305 VSS.n1157 VSS.t151 955.091
R2306 VSS.n1139 VSS.t223 955.091
R2307 VSS.n1146 VSS.t529 955.091
R2308 VSS.n1128 VSS.t416 955.091
R2309 VSS.n1135 VSS.t164 955.091
R2310 VSS.n1117 VSS.t177 955.091
R2311 VSS.n1124 VSS.t472 955.091
R2312 VSS.n1106 VSS.t411 955.091
R2313 VSS.n1113 VSS.t345 955.091
R2314 VSS.n1095 VSS.t484 955.091
R2315 VSS.n1102 VSS.t383 955.091
R2316 VSS.n805 VSS.t241 955.091
R2317 VSS.t441 VSS.n726 955.091
R2318 VSS.n1162 VSS.t195 935.33
R2319 VSS.n1151 VSS.t258 935.33
R2320 VSS.n1140 VSS.t494 935.33
R2321 VSS.n1129 VSS.t116 935.33
R2322 VSS.n1118 VSS.t29 935.33
R2323 VSS.n1107 VSS.t147 935.33
R2324 VSS.n1096 VSS.t118 935.33
R2325 VSS.n806 VSS.t375 935.33
R2326 VSS.n1091 VSS.n727 832.486
R2327 VSS.n873 VSS.n711 832.486
R2328 VSS.n1069 VSS.n696 832.486
R2329 VSS.n1035 VSS.n681 832.486
R2330 VSS.n991 VSS.n666 832.486
R2331 VSS.n957 VSS.n651 832.486
R2332 VSS.n913 VSS.n636 832.486
R2333 VSS.n1197 VSS.t189 815.229
R2334 VSS.n110 VSS.t496 815.229
R2335 VSS.t354 VSS.n110 815.229
R2336 VSS.n1200 VSS.t70 815.229
R2337 VSS.n945 VSS.t63 815.229
R2338 VSS.t556 VSS.n943 815.229
R2339 VSS.n943 VSS.t253 815.229
R2340 VSS.n1215 VSS.t460 815.229
R2341 VSS.n940 VSS.t464 815.229
R2342 VSS.t409 VSS.n940 815.229
R2343 VSS.n942 VSS.t391 815.229
R2344 VSS.n1218 VSS.t430 815.229
R2345 VSS.n1023 VSS.t511 815.229
R2346 VSS.t397 VSS.n1021 815.229
R2347 VSS.n1021 VSS.t288 815.229
R2348 VSS.n1233 VSS.t489 815.229
R2349 VSS.n1018 VSS.t373 815.229
R2350 VSS.t82 VSS.n1018 815.229
R2351 VSS.n1020 VSS.t294 815.229
R2352 VSS.n1236 VSS.t543 815.229
R2353 VSS.n749 VSS.t98 815.229
R2354 VSS.t68 VSS.n747 815.229
R2355 VSS.n747 VSS.t330 815.229
R2356 VSS.t311 VSS.n746 815.229
R2357 VSS.n764 VSS.t250 815.229
R2358 VSS.t335 VSS.n764 815.229
R2359 VSS.n765 VSS.t367 815.229
R2360 VSS.n112 VSS.t282 815.229
R2361 VSS.n632 VSS.t239 815.229
R2362 VSS.t560 VSS.n629 815.229
R2363 VSS.n629 VSS.t478 815.229
R2364 VSS.n521 VSS.n520 760.639
R2365 VSS.n524 VSS.n523 760.639
R2366 VSS.n550 VSS.n527 760.639
R2367 VSS.n564 VSS.n477 760.639
R2368 VSS.n559 VSS.n482 760.639
R2369 VSS.n485 VSS.n483 760.639
R2370 VSS.n488 VSS.n487 760.639
R2371 VSS.n308 VSS.n294 760.639
R2372 VSS.n312 VSS.n293 760.639
R2373 VSS.n321 VSS.n287 760.639
R2374 VSS.n325 VSS.n286 760.639
R2375 VSS.n334 VSS.n280 760.639
R2376 VSS.n338 VSS.n279 760.639
R2377 VSS.n347 VSS.n273 760.639
R2378 VSS.n351 VSS.n272 760.639
R2379 VSS.n360 VSS.n266 760.639
R2380 VSS.n364 VSS.n265 760.639
R2381 VSS.n373 VSS.n259 760.639
R2382 VSS.n377 VSS.n258 760.639
R2383 VSS.n386 VSS.n252 760.639
R2384 VSS.n390 VSS.n251 760.639
R2385 VSS.n399 VSS.n245 760.639
R2386 VSS.n403 VSS.n244 760.639
R2387 VSS.n412 VSS.n238 760.639
R2388 VSS.n416 VSS.n237 760.639
R2389 VSS.n425 VSS.n231 760.639
R2390 VSS.n429 VSS.n230 760.639
R2391 VSS.n438 VSS.n224 760.639
R2392 VSS.n442 VSS.n223 760.639
R2393 VSS.n451 VSS.n217 760.639
R2394 VSS.n455 VSS.n216 760.639
R2395 VSS.n466 VSS.n210 760.639
R2396 VSS.n470 VSS.n209 760.639
R2397 VSS.n475 VSS.n203 760.639
R2398 VSS.n911 VSS.n899 742.855
R2399 VSS.n955 VSS.n933 742.855
R2400 VSS.n989 VSS.n977 742.855
R2401 VSS.n1033 VSS.n1011 742.855
R2402 VSS.n1067 VSS.n1055 742.855
R2403 VSS.n864 VSS.n861 742.855
R2404 VSS.n104 VSS.n84 742.855
R2405 VSS.n834 VSS.n739 742.855
R2406 VSS.n619 VSS.n618 631.795
R2407 VSS.n152 VSS.n150 631.795
R2408 VSS.n603 VSS.n602 631.795
R2409 VSS.n178 VSS.n176 631.795
R2410 VSS.n587 VSS.n586 631.795
R2411 VSS.n515 VSS.n512 631.795
R2412 VSS.n1158 VSS.n1157 605.989
R2413 VSS.n1147 VSS.n1146 605.989
R2414 VSS.n1136 VSS.n1135 605.989
R2415 VSS.n1125 VSS.n1124 605.989
R2416 VSS.n1114 VSS.n1113 605.989
R2417 VSS.n1103 VSS.n1102 605.989
R2418 VSS.n1092 VSS.n726 605.989
R2419 VSS.n1159 VSS.n1158 592.814
R2420 VSS.n1148 VSS.n1147 592.814
R2421 VSS.n1137 VSS.n1136 592.814
R2422 VSS.n1126 VSS.n1125 592.814
R2423 VSS.n1115 VSS.n1114 592.814
R2424 VSS.n1104 VSS.n1103 592.814
R2425 VSS.n1093 VSS.n1092 592.814
R2426 VSS.t209 VSS.t262 579.641
R2427 VSS.t27 VSS.t209 579.641
R2428 VSS.t195 VSS.t27 579.641
R2429 VSS.t260 VSS.t493 579.641
R2430 VSS.t493 VSS.t280 579.641
R2431 VSS.t280 VSS.t371 579.641
R2432 VSS.t558 VSS.t343 579.641
R2433 VSS.t581 VSS.t558 579.641
R2434 VSS.t258 VSS.t581 579.641
R2435 VSS.t305 VSS.t107 579.641
R2436 VSS.t107 VSS.t7 579.641
R2437 VSS.t7 VSS.t151 579.641
R2438 VSS.t278 VSS.t419 579.641
R2439 VSS.t521 VSS.t278 579.641
R2440 VSS.t494 VSS.t521 579.641
R2441 VSS.t223 VSS.t536 579.641
R2442 VSS.t536 VSS.t172 579.641
R2443 VSS.t172 VSS.t529 579.641
R2444 VSS.t243 VSS.t0 579.641
R2445 VSS.t161 VSS.t243 579.641
R2446 VSS.t116 VSS.t161 579.641
R2447 VSS.t416 VSS.t3 579.641
R2448 VSS.t3 VSS.t270 579.641
R2449 VSS.t270 VSS.t164 579.641
R2450 VSS.t553 VSS.t470 579.641
R2451 VSS.t468 VSS.t553 579.641
R2452 VSS.t29 VSS.t468 579.641
R2453 VSS.t177 VSS.t469 579.641
R2454 VSS.t469 VSS.t482 579.641
R2455 VSS.t482 VSS.t472 579.641
R2456 VSS.t509 VSS.t112 579.641
R2457 VSS.t418 VSS.t509 579.641
R2458 VSS.t147 VSS.t418 579.641
R2459 VSS.t411 VSS.t351 579.641
R2460 VSS.t351 VSS.t124 579.641
R2461 VSS.t124 VSS.t345 579.641
R2462 VSS.t14 VSS.t387 579.641
R2463 VSS.t381 VSS.t14 579.641
R2464 VSS.t118 VSS.t381 579.641
R2465 VSS.t484 VSS.t386 579.641
R2466 VSS.t386 VSS.t389 579.641
R2467 VSS.t389 VSS.t383 579.641
R2468 VSS.t564 VSS.t378 579.641
R2469 VSS.t578 VSS.t564 579.641
R2470 VSS.t375 VSS.t578 579.641
R2471 VSS.t241 VSS.t380 579.641
R2472 VSS.t380 VSS.t225 579.641
R2473 VSS.t225 VSS.t441 579.641
R2474 VSS.n127 VSS.t166 549.061
R2475 VSS.t426 VSS.n127 549.061
R2476 VSS.n619 VSS.t534 549.061
R2477 VSS.n618 VSS.t369 549.061
R2478 VSS.n148 VSS.t214 549.061
R2479 VSS.t114 VSS.n148 549.061
R2480 VSS.n150 VSS.t434 549.061
R2481 VSS.t405 VSS.n152 549.061
R2482 VSS.n153 VSS.t54 549.061
R2483 VSS.t532 VSS.n153 549.061
R2484 VSS.n603 VSS.t100 549.061
R2485 VSS.n602 VSS.t357 549.061
R2486 VSS.n174 VSS.t105 549.061
R2487 VSS.t401 VSS.n174 549.061
R2488 VSS.n176 VSS.t136 549.061
R2489 VSS.t153 VSS.n178 549.061
R2490 VSS.n179 VSS.t579 549.061
R2491 VSS.t513 VSS.n179 549.061
R2492 VSS.n587 VSS.t315 549.061
R2493 VSS.n586 VSS.t140 549.061
R2494 VSS.n510 VSS.t48 549.061
R2495 VSS.t476 VSS.n510 549.061
R2496 VSS.n512 VSS.t91 549.061
R2497 VSS.t571 VSS.n515 549.061
R2498 VSS.n516 VSS.t451 549.061
R2499 VSS.t193 VSS.n516 549.061
R2500 VSS.n827 VSS.n826 546.538
R2501 VSS.n509 VSS.n508 509.743
R2502 VSS.t525 VSS.t189 491.372
R2503 VSS.t159 VSS.t525 491.372
R2504 VSS.t496 VSS.t159 491.372
R2505 VSS.t181 VSS.t421 491.372
R2506 VSS.t421 VSS.t70 491.372
R2507 VSS.t63 VSS.t87 491.372
R2508 VSS.t87 VSS.t569 491.372
R2509 VSS.t569 VSS.t556 491.372
R2510 VSS.t466 VSS.t460 491.372
R2511 VSS.t458 VSS.t466 491.372
R2512 VSS.t464 VSS.t458 491.372
R2513 VSS.t407 VSS.t567 491.372
R2514 VSS.t391 VSS.t407 491.372
R2515 VSS.t573 VSS.t576 491.372
R2516 VSS.t576 VSS.t430 491.372
R2517 VSS.t511 VSS.t395 491.372
R2518 VSS.t395 VSS.t393 491.372
R2519 VSS.t393 VSS.t397 491.372
R2520 VSS.t297 VSS.t489 491.372
R2521 VSS.t149 VSS.t297 491.372
R2522 VSS.t373 VSS.t149 491.372
R2523 VSS.t145 VSS.t79 491.372
R2524 VSS.t294 VSS.t145 491.372
R2525 VSS.t541 VSS.t328 491.372
R2526 VSS.t328 VSS.t543 491.372
R2527 VSS.t98 VSS.t51 491.372
R2528 VSS.t51 VSS.t403 491.372
R2529 VSS.t403 VSS.t68 491.372
R2530 VSS.t453 VSS.t311 491.372
R2531 VSS.t456 VSS.t453 491.372
R2532 VSS.t250 VSS.t456 491.372
R2533 VSS.t268 VSS.t127 491.372
R2534 VSS.t367 VSS.t268 491.372
R2535 VSS.t486 VSS.t491 491.372
R2536 VSS.t282 VSS.t486 491.372
R2537 VSS.t239 VSS.t264 491.372
R2538 VSS.t264 VSS.t217 491.372
R2539 VSS.t217 VSS.t560 491.372
R2540 VSS.t491 VSS.t354 477.411
R2541 VSS.t253 VSS.t181 477.411
R2542 VSS.t567 VSS.t409 477.411
R2543 VSS.t288 VSS.t573 477.411
R2544 VSS.t79 VSS.t82 477.411
R2545 VSS.t330 VSS.t541 477.411
R2546 VSS.t127 VSS.t335 477.411
R2547 VSS.t478 VSS.t272 471.786
R2548 VSS.n1090 VSS.n1089 446.182
R2549 VSS.n1062 VSS.n11 446.182
R2550 VSS.n1028 VSS.n1027 446.182
R2551 VSS.n984 VSS.n33 446.182
R2552 VSS.n950 VSS.n949 446.182
R2553 VSS.n906 VSS.n55 446.182
R2554 VSS.n635 VSS.n109 446.182
R2555 VSS.n1091 VSS.n1090 413.346
R2556 VSS.n711 VSS.n11 413.346
R2557 VSS.n1027 VSS.n696 413.346
R2558 VSS.n681 VSS.n33 413.346
R2559 VSS.n949 VSS.n666 413.346
R2560 VSS.n651 VSS.n55 413.346
R2561 VSS.n636 VSS.n635 413.346
R2562 VSS.n908 VSS.n899 356.277
R2563 VSS.n952 VSS.n933 356.277
R2564 VSS.n986 VSS.n977 356.277
R2565 VSS.n1030 VSS.n1011 356.277
R2566 VSS.n1064 VSS.n1055 356.277
R2567 VSS.n861 VSS.n729 356.277
R2568 VSS.n107 VSS.n84 356.277
R2569 VSS.n830 VSS.n739 356.277
R2570 VSS.t256 VSS.n628 346.868
R2571 VSS.n625 VSS.t155 346.868
R2572 VSS.t41 VSS.n727 338.017
R2573 VSS.n1089 VSS.t303 338.017
R2574 VSS.n873 VSS.t382 338.017
R2575 VSS.t170 VSS.n1062 338.017
R2576 VSS.t235 VSS.n1069 338.017
R2577 VSS.t212 VSS.n1028 338.017
R2578 VSS.t42 VSS.n1035 338.017
R2579 VSS.t207 VSS.n984 338.017
R2580 VSS.t162 VSS.n991 338.017
R2581 VSS.t33 VSS.n950 338.017
R2582 VSS.t102 VSS.n957 338.017
R2583 VSS.t76 VSS.n906 338.017
R2584 VSS.t555 VSS.n913 338.017
R2585 VSS.n109 VSS.t266 338.017
R2586 VSS.t166 VSS.t157 330.94
R2587 VSS.t474 VSS.t426 330.94
R2588 VSS.t191 VSS.t474 330.94
R2589 VSS.t534 VSS.t191 330.94
R2590 VSS.t24 VSS.t369 330.94
R2591 VSS.t505 VSS.t24 330.94
R2592 VSS.t214 VSS.t505 330.94
R2593 VSS.t349 VSS.t114 330.94
R2594 VSS.t436 VSS.t349 330.94
R2595 VSS.t434 VSS.t436 330.94
R2596 VSS.t547 VSS.t405 330.94
R2597 VSS.t549 VSS.t547 330.94
R2598 VSS.t54 VSS.t549 330.94
R2599 VSS.t286 VSS.t532 330.94
R2600 VSS.t399 VSS.t286 330.94
R2601 VSS.t100 VSS.t399 330.94
R2602 VSS.t447 VSS.t357 330.94
R2603 VSS.t284 VSS.t447 330.94
R2604 VSS.t105 VSS.t284 330.94
R2605 VSS.t449 VSS.t401 330.94
R2606 VSS.t527 VSS.t449 330.94
R2607 VSS.t136 VSS.t527 330.94
R2608 VSS.t562 VSS.t153 330.94
R2609 VSS.t582 VSS.t562 330.94
R2610 VSS.t579 VSS.t582 330.94
R2611 VSS.t507 VSS.t513 330.94
R2612 VSS.t428 VSS.t507 330.94
R2613 VSS.t315 VSS.t428 330.94
R2614 VSS.t175 VSS.t140 330.94
R2615 VSS.t93 VSS.t175 330.94
R2616 VSS.t48 VSS.t93 330.94
R2617 VSS.t290 VSS.t476 330.94
R2618 VSS.t66 VSS.t290 330.94
R2619 VSS.t91 VSS.t66 330.94
R2620 VSS.t39 VSS.t571 330.94
R2621 VSS.t309 VSS.t39 330.94
R2622 VSS.t451 VSS.t309 330.94
R2623 VSS.t499 VSS.t193 330.94
R2624 VSS.n517 VSS.t89 317.079
R2625 VSS.t424 VSS.n518 314.906
R2626 VSS.n565 VSS.t18 314.906
R2627 VSS.n521 VSS.n519 297.553
R2628 VSS.n522 VSS.n521 297.553
R2629 VSS.n524 VSS.n522 297.553
R2630 VSS.n525 VSS.n524 297.553
R2631 VSS.n527 VSS.n525 297.553
R2632 VSS.n527 VSS.n526 297.553
R2633 VSS.n526 VSS.n477 297.553
R2634 VSS.n560 VSS.n477 297.553
R2635 VSS.n560 VSS.n559 297.553
R2636 VSS.n559 VSS.n558 297.553
R2637 VSS.n558 VSS.n483 297.553
R2638 VSS.n486 VSS.n483 297.553
R2639 VSS.n488 VSS.n486 297.553
R2640 VSS.n489 VSS.n488 297.553
R2641 VSS.n300 VSS.n294 297.553
R2642 VSS.n311 VSS.n294 297.553
R2643 VSS.n312 VSS.n311 297.553
R2644 VSS.n313 VSS.n312 297.553
R2645 VSS.n313 VSS.n287 297.553
R2646 VSS.n324 VSS.n287 297.553
R2647 VSS.n325 VSS.n324 297.553
R2648 VSS.n326 VSS.n325 297.553
R2649 VSS.n326 VSS.n280 297.553
R2650 VSS.n337 VSS.n280 297.553
R2651 VSS.n338 VSS.n337 297.553
R2652 VSS.n339 VSS.n338 297.553
R2653 VSS.n339 VSS.n273 297.553
R2654 VSS.n350 VSS.n273 297.553
R2655 VSS.n351 VSS.n350 297.553
R2656 VSS.n352 VSS.n351 297.553
R2657 VSS.n352 VSS.n266 297.553
R2658 VSS.n363 VSS.n266 297.553
R2659 VSS.n364 VSS.n363 297.553
R2660 VSS.n365 VSS.n364 297.553
R2661 VSS.n365 VSS.n259 297.553
R2662 VSS.n376 VSS.n259 297.553
R2663 VSS.n377 VSS.n376 297.553
R2664 VSS.n378 VSS.n377 297.553
R2665 VSS.n378 VSS.n252 297.553
R2666 VSS.n389 VSS.n252 297.553
R2667 VSS.n390 VSS.n389 297.553
R2668 VSS.n391 VSS.n390 297.553
R2669 VSS.n391 VSS.n245 297.553
R2670 VSS.n402 VSS.n245 297.553
R2671 VSS.n403 VSS.n402 297.553
R2672 VSS.n404 VSS.n403 297.553
R2673 VSS.n404 VSS.n238 297.553
R2674 VSS.n415 VSS.n238 297.553
R2675 VSS.n416 VSS.n415 297.553
R2676 VSS.n417 VSS.n416 297.553
R2677 VSS.n417 VSS.n231 297.553
R2678 VSS.n428 VSS.n231 297.553
R2679 VSS.n429 VSS.n428 297.553
R2680 VSS.n430 VSS.n429 297.553
R2681 VSS.n430 VSS.n224 297.553
R2682 VSS.n441 VSS.n224 297.553
R2683 VSS.n442 VSS.n441 297.553
R2684 VSS.n443 VSS.n442 297.553
R2685 VSS.n443 VSS.n217 297.553
R2686 VSS.n454 VSS.n217 297.553
R2687 VSS.n455 VSS.n454 297.553
R2688 VSS.n456 VSS.n455 297.553
R2689 VSS.n456 VSS.n210 297.553
R2690 VSS.n469 VSS.n210 297.553
R2691 VSS.n470 VSS.n469 297.553
R2692 VSS.n471 VSS.n470 297.553
R2693 VSS.n471 VSS.n203 297.553
R2694 VSS.n203 VSS.n202 297.553
R2695 VSS.n832 VSS.n746 295.94
R2696 VSS.n553 VSS.t432 291.325
R2697 VSS.n552 VSS.t438 291.325
R2698 VSS.n551 VSS.t16 291.325
R2699 VSS.t20 VSS.n556 291.325
R2700 VSS.t22 VSS.n555 291.325
R2701 VSS.t424 VSS.n553 291.325
R2702 VSS.t432 VSS.n552 291.325
R2703 VSS.t438 VSS.n551 291.325
R2704 VSS.t20 VSS.n557 291.325
R2705 VSS.n556 VSS.t22 291.325
R2706 VSS.n555 VSS.t537 291.325
R2707 VSS.n557 VSS.t18 291.325
R2708 VSS.n904 VSS.n897 281.135
R2709 VSS.n938 VSS.n931 281.135
R2710 VSS.n982 VSS.n975 281.135
R2711 VSS.n1016 VSS.n1009 281.135
R2712 VSS.n1060 VSS.n1053 281.135
R2713 VSS.n874 VSS.n855 281.135
R2714 VSS.n89 VSS.n82 281.135
R2715 VSS.n744 VSS.n737 281.135
R2716 VSS.t322 VSS.t499 275.329
R2717 VSS.n743 VSS.n742 262.659
R2718 VSS.n859 VSS.n854 262.659
R2719 VSS.n1059 VSS.n1058 262.659
R2720 VSS.n1015 VSS.n1014 262.659
R2721 VSS.n981 VSS.n980 262.659
R2722 VSS.n937 VSS.n936 262.659
R2723 VSS.n903 VSS.n902 262.659
R2724 VSS.n88 VSS.n87 262.659
R2725 VSS.t157 VSS.t443 246.464
R2726 VSS.t28 VSS.n1170 218.262
R2727 VSS.n566 VSS.t16 217.178
R2728 VSS.t272 VSS.t103 209.071
R2729 VSS.t103 VSS.t256 209.071
R2730 VSS.t443 VSS.t155 209.071
R2731 VSS.n553 VSS.n520 206.792
R2732 VSS.n552 VSS.n523 206.792
R2733 VSS.n551 VSS.n550 206.792
R2734 VSS.n556 VSS.n485 206.792
R2735 VSS.n555 VSS.n487 206.792
R2736 VSS.n557 VSS.n482 206.71
R2737 VSS.n745 VSS.n743 204.031
R2738 VSS.n863 VSS.n859 204.031
R2739 VSS.n1061 VSS.n1059 204.031
R2740 VSS.n1017 VSS.n1015 204.031
R2741 VSS.n983 VSS.n981 204.031
R2742 VSS.n939 VSS.n937 204.031
R2743 VSS.n905 VSS.n903 204.031
R2744 VSS.n103 VSS.n88 204.031
R2745 VSS.n844 VSS.n732 202.725
R2746 VSS.n1086 VSS.n1085 202.725
R2747 VSS.n1078 VSS.n1051 202.725
R2748 VSS.n1044 VSS.n1007 202.725
R2749 VSS.n1000 VSS.n973 202.725
R2750 VSS.n966 VSS.n929 202.725
R2751 VSS.n922 VSS.n895 202.725
R2752 VSS.n1179 VSS.n77 202.725
R2753 VSS.n475 VSS.n474 195
R2754 VSS.n476 VSS.n475 195
R2755 VSS.n460 VSS.n209 195
R2756 VSS.n468 VSS.n209 195
R2757 VSS.n466 VSS.n465 195
R2758 VSS.n467 VSS.n466 195
R2759 VSS.n216 VSS.n215 195
R2760 VSS.n453 VSS.n216 195
R2761 VSS.n451 VSS.n450 195
R2762 VSS.n452 VSS.n451 195
R2763 VSS.n223 VSS.n222 195
R2764 VSS.n440 VSS.n223 195
R2765 VSS.n438 VSS.n437 195
R2766 VSS.n439 VSS.n438 195
R2767 VSS.n230 VSS.n229 195
R2768 VSS.n427 VSS.n230 195
R2769 VSS.n425 VSS.n424 195
R2770 VSS.n426 VSS.n425 195
R2771 VSS.n237 VSS.n236 195
R2772 VSS.n414 VSS.n237 195
R2773 VSS.n412 VSS.n411 195
R2774 VSS.n413 VSS.n412 195
R2775 VSS.n244 VSS.n243 195
R2776 VSS.n401 VSS.n244 195
R2777 VSS.n399 VSS.n398 195
R2778 VSS.n400 VSS.n399 195
R2779 VSS.n251 VSS.n250 195
R2780 VSS.n388 VSS.n251 195
R2781 VSS.n386 VSS.n385 195
R2782 VSS.n387 VSS.n386 195
R2783 VSS.n258 VSS.n257 195
R2784 VSS.n375 VSS.n258 195
R2785 VSS.n373 VSS.n372 195
R2786 VSS.n374 VSS.n373 195
R2787 VSS.n265 VSS.n264 195
R2788 VSS.n362 VSS.n265 195
R2789 VSS.n360 VSS.n359 195
R2790 VSS.n361 VSS.n360 195
R2791 VSS.n272 VSS.n271 195
R2792 VSS.n349 VSS.n272 195
R2793 VSS.n347 VSS.n346 195
R2794 VSS.n348 VSS.n347 195
R2795 VSS.n279 VSS.n278 195
R2796 VSS.n336 VSS.n279 195
R2797 VSS.n334 VSS.n333 195
R2798 VSS.n335 VSS.n334 195
R2799 VSS.n286 VSS.n285 195
R2800 VSS.n323 VSS.n286 195
R2801 VSS.n321 VSS.n320 195
R2802 VSS.n322 VSS.n321 195
R2803 VSS.n293 VSS.n292 195
R2804 VSS.n310 VSS.n293 195
R2805 VSS.n308 VSS.n307 195
R2806 VSS.n309 VSS.n308 195
R2807 VSS.n299 VSS.n298 195
R2808 VSS.n299 VSS.n92 195
R2809 VSS.n569 VSS.n568 195
R2810 VSS.n568 VSS.n567 195
R2811 VSS.n491 VSS.n487 195
R2812 VSS.n498 VSS.n485 195
R2813 VSS.n492 VSS.n482 195
R2814 VSS.n564 VSS.n563 195
R2815 VSS.n565 VSS.n564 195
R2816 VSS.n550 VSS.n549 195
R2817 VSS.n532 VSS.n523 195
R2818 VSS.n534 VSS.n520 195
R2819 VSS.n536 VSS.n535 195
R2820 VSS.n535 VSS.n518 195
R2821 VSS.t89 VSS.t322 191.115
R2822 VSS.t168 VSS.n828 186.441
R2823 VSS.t501 VSS.n92 170.954
R2824 VSS.n309 VSS.t501 170.954
R2825 VSS.t95 VSS.n309 170.954
R2826 VSS.t95 VSS.n310 170.954
R2827 VSS.n310 VSS.t197 170.954
R2828 VSS.n322 VSS.t197 170.954
R2829 VSS.t519 VSS.n322 170.954
R2830 VSS.t519 VSS.n323 170.954
R2831 VSS.n323 VSS.t539 170.954
R2832 VSS.n335 VSS.t539 170.954
R2833 VSS.t221 VSS.n335 170.954
R2834 VSS.t221 VSS.n336 170.954
R2835 VSS.n336 VSS.t361 170.954
R2836 VSS.n348 VSS.t361 170.954
R2837 VSS.t326 VSS.n348 170.954
R2838 VSS.t326 VSS.n349 170.954
R2839 VSS.n349 VSS.t122 170.954
R2840 VSS.n361 VSS.t122 170.954
R2841 VSS.t5 VSS.n361 170.954
R2842 VSS.t5 VSS.n362 170.954
R2843 VSS.n362 VSS.t43 170.954
R2844 VSS.n374 VSS.t43 170.954
R2845 VSS.t120 VSS.n374 170.954
R2846 VSS.t120 VSS.n375 170.954
R2847 VSS.n375 VSS.t324 170.954
R2848 VSS.n387 VSS.t324 170.954
R2849 VSS.t517 VSS.n387 170.954
R2850 VSS.t517 VSS.n388 170.954
R2851 VSS.n388 VSS.t199 170.954
R2852 VSS.n400 VSS.t199 170.954
R2853 VSS.t219 VSS.n400 170.954
R2854 VSS.t219 VSS.n401 170.954
R2855 VSS.n401 VSS.t229 170.954
R2856 VSS.n413 VSS.t229 170.954
R2857 VSS.t233 VSS.n413 170.954
R2858 VSS.t233 VSS.n414 170.954
R2859 VSS.n414 VSS.t231 170.954
R2860 VSS.n426 VSS.t231 170.954
R2861 VSS.t227 VSS.n426 170.954
R2862 VSS.t227 VSS.n427 170.954
R2863 VSS.n427 VSS.t58 170.954
R2864 VSS.n439 VSS.t58 170.954
R2865 VSS.t10 VSS.n439 170.954
R2866 VSS.t10 VSS.n440 170.954
R2867 VSS.n440 VSS.t183 170.954
R2868 VSS.n452 VSS.t183 170.954
R2869 VSS.t274 VSS.n452 170.954
R2870 VSS.t274 VSS.n453 170.954
R2871 VSS.n453 VSS.t143 170.954
R2872 VSS.n467 VSS.t143 170.954
R2873 VSS.t313 VSS.n467 170.954
R2874 VSS.t313 VSS.n468 170.954
R2875 VSS.n468 VSS.t445 170.954
R2876 VSS.n476 VSS.t445 170.954
R2877 VSS.t515 VSS.n476 170.954
R2878 VSS.n567 VSS.t515 170.954
R2879 VSS.t413 VSS.t35 169.975
R2880 VSS.t35 VSS.t47 169.975
R2881 VSS.t377 VSS.t47 169.975
R2882 VSS.t377 VSS.t423 169.975
R2883 VSS.t423 VSS.t131 169.975
R2884 VSS.t75 VSS.t206 169.975
R2885 VSS.t206 VSS.t440 169.975
R2886 VSS.t440 VSS.t41 169.975
R2887 VSS.t31 VSS.t84 169.975
R2888 VSS.t503 VSS.t12 169.975
R2889 VSS.t385 VSS.t503 169.975
R2890 VSS.t216 VSS.t385 169.975
R2891 VSS.t72 VSS.t216 169.975
R2892 VSS.t455 VSS.t72 169.975
R2893 VSS.t126 VSS.t334 169.975
R2894 VSS.t252 VSS.t126 169.975
R2895 VSS.t382 VSS.t252 169.975
R2896 VSS.t202 VSS.t237 169.975
R2897 VSS.t134 VSS.t480 169.975
R2898 VSS.t480 VSS.t321 169.975
R2899 VSS.t174 VSS.t321 169.975
R2900 VSS.t174 VSS.t142 169.975
R2901 VSS.t142 VSS.t97 169.975
R2902 VSS.t53 VSS.t201 169.975
R2903 VSS.t201 VSS.t50 169.975
R2904 VSS.t50 VSS.t235 169.975
R2905 VSS.t187 VSS.t359 169.975
R2906 VSS.t301 VSS.t245 169.975
R2907 VSS.t245 VSS.t81 169.975
R2908 VSS.t78 VSS.t81 169.975
R2909 VSS.t78 VSS.t522 169.975
R2910 VSS.t522 VSS.t300 169.975
R2911 VSS.t60 VSS.t415 169.975
R2912 VSS.t415 VSS.t108 169.975
R2913 VSS.t108 VSS.t42 169.975
R2914 VSS.t37 VSS.t551 169.975
R2915 VSS.t185 VSS.t247 169.975
R2916 VSS.t247 VSS.t4 169.975
R2917 VSS.t2 VSS.t4 169.975
R2918 VSS.t2 VSS.t523 169.975
R2919 VSS.t523 VSS.t524 169.975
R2920 VSS.t488 VSS.t575 169.975
R2921 VSS.t575 VSS.t163 169.975
R2922 VSS.t163 VSS.t162 169.975
R2923 VSS.t545 VSS.t363 169.975
R2924 VSS.t347 VSS.t276 169.975
R2925 VSS.t276 VSS.t26 169.975
R2926 VSS.t255 VSS.t26 169.975
R2927 VSS.t255 VSS.t462 169.975
R2928 VSS.t462 VSS.t463 169.975
R2929 VSS.t566 VSS.t9 169.975
R2930 VSS.t9 VSS.t111 169.975
R2931 VSS.t111 VSS.t102 169.975
R2932 VSS.t332 VSS.t132 169.975
R2933 VSS.t73 VSS.t341 169.975
R2934 VSS.t341 VSS.t299 169.975
R2935 VSS.t110 VSS.t299 169.975
R2936 VSS.t110 VSS.t211 169.975
R2937 VSS.t211 VSS.t65 169.975
R2938 VSS.t236 VSS.t109 169.975
R2939 VSS.t109 VSS.t86 169.975
R2940 VSS.t86 VSS.t555 169.975
R2941 VSS.t292 VSS.t352 169.975
R2942 VSS.t337 VSS.t56 169.975
R2943 VSS.t56 VSS.t307 169.975
R2944 VSS.t308 VSS.t307 169.975
R2945 VSS.t308 VSS.t531 169.975
R2946 VSS.t531 VSS.t356 169.975
R2947 VSS.t498 VSS.t249 169.975
R2948 VSS.t249 VSS.t296 169.975
R2949 VSS.t296 VSS.t28 169.975
R2950 VSS.n865 VSS.t31 168.042
R2951 VSS.n1066 VSS.t202 168.042
R2952 VSS.n1032 VSS.t187 168.042
R2953 VSS.n988 VSS.t37 168.042
R2954 VSS.n954 VSS.t545 168.042
R2955 VSS.n910 VSS.t332 168.042
R2956 VSS.t352 VSS.n105 168.042
R2957 VSS.t319 VSS.n799 155.546
R2958 VSS.n800 VSS.t61 155.546
R2959 VSS.n826 VSS.t204 155.546
R2960 VSS.n844 VSS.n735 152.744
R2961 VSS.n1087 VSS.n1086 152.744
R2962 VSS.n1078 VSS.n875 152.744
R2963 VSS.n1044 VSS.n878 152.744
R2964 VSS.n1000 VSS.n881 152.744
R2965 VSS.n966 VSS.n884 152.744
R2966 VSS.n922 VSS.n887 152.744
R2967 VSS.n1179 VSS.n80 152.744
R2968 VSS.n621 VSS.n620 146.25
R2969 VSS.n620 VSS.n619 146.25
R2970 VSS.n617 VSS.n616 146.25
R2971 VSS.n618 VSS.n617 146.25
R2972 VSS.n149 VSS.n131 146.25
R2973 VSS.n150 VSS.n149 146.25
R2974 VSS.n151 VSS.n138 146.25
R2975 VSS.n152 VSS.n151 146.25
R2976 VSS.n605 VSS.n604 146.25
R2977 VSS.n604 VSS.n603 146.25
R2978 VSS.n601 VSS.n600 146.25
R2979 VSS.n602 VSS.n601 146.25
R2980 VSS.n175 VSS.n157 146.25
R2981 VSS.n176 VSS.n175 146.25
R2982 VSS.n177 VSS.n164 146.25
R2983 VSS.n178 VSS.n177 146.25
R2984 VSS.n589 VSS.n588 146.25
R2985 VSS.n588 VSS.n587 146.25
R2986 VSS.n585 VSS.n584 146.25
R2987 VSS.n586 VSS.n585 146.25
R2988 VSS.n511 VSS.n183 146.25
R2989 VSS.n512 VSS.n511 146.25
R2990 VSS.n514 VSS.n190 146.25
R2991 VSS.n515 VSS.n514 146.25
R2992 VSS.n1196 VSS.n1195 146.25
R2993 VSS.n1197 VSS.n1196 146.25
R2994 VSS.n1202 VSS.n1201 146.25
R2995 VSS.n1201 VSS.n1200 146.25
R2996 VSS.n944 VSS.n45 146.25
R2997 VSS.n945 VSS.n944 146.25
R2998 VSS.n1214 VSS.n1213 146.25
R2999 VSS.n1215 VSS.n1214 146.25
R3000 VSS.n941 VSS.n38 146.25
R3001 VSS.n942 VSS.n941 146.25
R3002 VSS.n1220 VSS.n1219 146.25
R3003 VSS.n1219 VSS.n1218 146.25
R3004 VSS.n1022 VSS.n23 146.25
R3005 VSS.n1023 VSS.n1022 146.25
R3006 VSS.n1232 VSS.n1231 146.25
R3007 VSS.n1233 VSS.n1232 146.25
R3008 VSS.n1019 VSS.n16 146.25
R3009 VSS.n1020 VSS.n1019 146.25
R3010 VSS.n1238 VSS.n1237 146.25
R3011 VSS.n1237 VSS.n1236 146.25
R3012 VSS.n748 VSS.n1 146.25
R3013 VSS.n749 VSS.n748 146.25
R3014 VSS.n762 VSS.n754 146.25
R3015 VSS.n762 VSS.n746 146.25
R3016 VSS.n767 VSS.n766 146.25
R3017 VSS.n766 VSS.n765 146.25
R3018 VSS.n798 VSS.n775 146.25
R3019 VSS.n799 VSS.n798 146.25
R3020 VSS.n825 VSS.n824 146.25
R3021 VSS.n826 VSS.n825 146.25
R3022 VSS.n301 VSS.n300 146.25
R3023 VSS.n300 VSS.t501 146.25
R3024 VSS.n311 VSS.n295 146.25
R3025 VSS.n311 VSS.t95 146.25
R3026 VSS.n314 VSS.n313 146.25
R3027 VSS.n313 VSS.t197 146.25
R3028 VSS.n324 VSS.n288 146.25
R3029 VSS.n324 VSS.t519 146.25
R3030 VSS.n327 VSS.n326 146.25
R3031 VSS.n326 VSS.t539 146.25
R3032 VSS.n337 VSS.n281 146.25
R3033 VSS.n337 VSS.t221 146.25
R3034 VSS.n340 VSS.n339 146.25
R3035 VSS.n339 VSS.t361 146.25
R3036 VSS.n350 VSS.n274 146.25
R3037 VSS.n350 VSS.t326 146.25
R3038 VSS.n353 VSS.n352 146.25
R3039 VSS.n352 VSS.t122 146.25
R3040 VSS.n363 VSS.n267 146.25
R3041 VSS.n363 VSS.t5 146.25
R3042 VSS.n366 VSS.n365 146.25
R3043 VSS.n365 VSS.t43 146.25
R3044 VSS.n376 VSS.n260 146.25
R3045 VSS.n376 VSS.t120 146.25
R3046 VSS.n379 VSS.n378 146.25
R3047 VSS.n378 VSS.t324 146.25
R3048 VSS.n389 VSS.n253 146.25
R3049 VSS.n389 VSS.t517 146.25
R3050 VSS.n392 VSS.n391 146.25
R3051 VSS.n391 VSS.t199 146.25
R3052 VSS.n402 VSS.n246 146.25
R3053 VSS.n402 VSS.t219 146.25
R3054 VSS.n405 VSS.n404 146.25
R3055 VSS.n404 VSS.t229 146.25
R3056 VSS.n415 VSS.n239 146.25
R3057 VSS.n415 VSS.t233 146.25
R3058 VSS.n418 VSS.n417 146.25
R3059 VSS.n417 VSS.t231 146.25
R3060 VSS.n428 VSS.n232 146.25
R3061 VSS.n428 VSS.t227 146.25
R3062 VSS.n431 VSS.n430 146.25
R3063 VSS.n430 VSS.t58 146.25
R3064 VSS.n441 VSS.n225 146.25
R3065 VSS.n441 VSS.t10 146.25
R3066 VSS.n444 VSS.n443 146.25
R3067 VSS.n443 VSS.t183 146.25
R3068 VSS.n454 VSS.n218 146.25
R3069 VSS.n454 VSS.t274 146.25
R3070 VSS.n457 VSS.n456 146.25
R3071 VSS.n456 VSS.t143 146.25
R3072 VSS.n469 VSS.n211 146.25
R3073 VSS.n469 VSS.t313 146.25
R3074 VSS.n472 VSS.n471 146.25
R3075 VSS.n471 VSS.t445 146.25
R3076 VSS.n202 VSS.n201 146.25
R3077 VSS.t515 VSS.n202 146.25
R3078 VSS.n573 VSS.n196 146.25
R3079 VSS.n517 VSS.n196 146.25
R3080 VSS.n539 VSS.n519 146.25
R3081 VSS.t424 VSS.n519 146.25
R3082 VSS.n541 VSS.n522 146.25
R3083 VSS.t432 VSS.n522 146.25
R3084 VSS.n547 VSS.n525 146.25
R3085 VSS.t438 VSS.n525 146.25
R3086 VSS.n526 VSS.n479 146.25
R3087 VSS.n526 VSS.t16 146.25
R3088 VSS.n561 VSS.n560 146.25
R3089 VSS.n560 VSS.t18 146.25
R3090 VSS.n558 VSS.n484 146.25
R3091 VSS.n558 VSS.t20 146.25
R3092 VSS.n501 VSS.n486 146.25
R3093 VSS.t22 VSS.n486 146.25
R3094 VSS.n490 VSS.n489 146.25
R3095 VSS.n624 VSS.n623 146.25
R3096 VSS.n625 VSS.n624 146.25
R3097 VSS.n111 VSS.n60 146.25
R3098 VSS.n112 VSS.n111 146.25
R3099 VSS.n631 VSS.n67 146.25
R3100 VSS.n632 VSS.n631 146.25
R3101 VSS.n1184 VSS.n73 146.25
R3102 VSS.n628 VSS.n73 146.25
R3103 VSS.n801 VSS.t339 142.761
R3104 VSS.n808 VSS.n782 136.387
R3105 VSS.n1098 VSS.n719 136.387
R3106 VSS.n1109 VSS.n704 136.387
R3107 VSS.n1120 VSS.n689 136.387
R3108 VSS.n1131 VSS.n674 136.387
R3109 VSS.n1142 VSS.n659 136.387
R3110 VSS.n1153 VSS.n644 136.387
R3111 VSS.n1164 VSS.n96 136.387
R3112 VSS.n795 VSS.n785 136.011
R3113 VSS.n1100 VSS.n1099 136.011
R3114 VSS.n1111 VSS.n1110 136.011
R3115 VSS.n1122 VSS.n1121 136.011
R3116 VSS.n1133 VSS.n1132 136.011
R3117 VSS.n1144 VSS.n1143 136.011
R3118 VSS.n1155 VSS.n1154 136.011
R3119 VSS.n1166 VSS.n1165 136.011
R3120 VSS.n583 VSS.n183 133.755
R3121 VSS.n584 VSS.n583 133.755
R3122 VSS.n590 VSS.n589 133.755
R3123 VSS.n590 VSS.n164 133.755
R3124 VSS.n599 VSS.n157 133.755
R3125 VSS.n600 VSS.n599 133.755
R3126 VSS.n606 VSS.n605 133.755
R3127 VSS.n606 VSS.n138 133.755
R3128 VSS.n615 VSS.n131 133.755
R3129 VSS.n616 VSS.n615 133.755
R3130 VSS.n623 VSS.n622 133.755
R3131 VSS.n622 VSS.n621 133.755
R3132 VSS.n574 VSS.n190 133.755
R3133 VSS.n574 VSS.n573 133.755
R3134 VSS.n824 VSS.n823 133.755
R3135 VSS.n823 VSS.n775 133.755
R3136 VSS.n1239 VSS.n1 133.755
R3137 VSS.n1239 VSS.n1238 133.755
R3138 VSS.n1221 VSS.n23 133.755
R3139 VSS.n1221 VSS.n1220 133.755
R3140 VSS.n1203 VSS.n45 133.755
R3141 VSS.n1203 VSS.n1202 133.755
R3142 VSS.n1194 VSS.n60 133.755
R3143 VSS.n1195 VSS.n1194 133.755
R3144 VSS.n1212 VSS.n38 133.755
R3145 VSS.n1213 VSS.n1212 133.755
R3146 VSS.n1230 VSS.n16 133.755
R3147 VSS.n1231 VSS.n1230 133.755
R3148 VSS.n768 VSS.n767 133.755
R3149 VSS.n768 VSS.n754 133.755
R3150 VSS.n1185 VSS.n67 133.755
R3151 VSS.n1185 VSS.n1184 133.755
R3152 VSS.n838 VSS.n743 124.481
R3153 VSS.n870 VSS.n859 124.481
R3154 VSS.n1072 VSS.n1059 124.481
R3155 VSS.n1038 VSS.n1015 124.481
R3156 VSS.n994 VSS.n981 124.481
R3157 VSS.n960 VSS.n937 124.481
R3158 VSS.n916 VSS.n903 124.481
R3159 VSS.n1173 VSS.n88 124.481
R3160 VSS.n839 VSS.n838 119.04
R3161 VSS.n870 VSS.n869 119.04
R3162 VSS.n1073 VSS.n1072 119.04
R3163 VSS.n1039 VSS.n1038 119.04
R3164 VSS.n995 VSS.n994 119.04
R3165 VSS.n961 VSS.n960 119.04
R3166 VSS.n917 VSS.n916 119.04
R3167 VSS.n1174 VSS.n1173 119.04
R3168 VSS.n830 VSS.n829 117.001
R3169 VSS.n831 VSS.n830 117.001
R3170 VSS.n731 VSS.n729 117.001
R3171 VSS.n862 VSS.n729 117.001
R3172 VSS.n1064 VSS.n1063 117.001
R3173 VSS.n1065 VSS.n1064 117.001
R3174 VSS.n1030 VSS.n1029 117.001
R3175 VSS.n1031 VSS.n1030 117.001
R3176 VSS.n986 VSS.n985 117.001
R3177 VSS.n987 VSS.n986 117.001
R3178 VSS.n952 VSS.n951 117.001
R3179 VSS.n953 VSS.n952 117.001
R3180 VSS.n908 VSS.n907 117.001
R3181 VSS.n909 VSS.n908 117.001
R3182 VSS.n107 VSS.n106 117.001
R3183 VSS.n108 VSS.n107 117.001
R3184 VSS.n627 VSS.n626 111.663
R3185 VSS.n829 VSS.n735 101.555
R3186 VSS.n1087 VSS.n731 101.555
R3187 VSS.n1063 VSS.n875 101.555
R3188 VSS.n1029 VSS.n878 101.555
R3189 VSS.n985 VSS.n881 101.555
R3190 VSS.n951 VSS.n884 101.555
R3191 VSS.n907 VSS.n887 101.555
R3192 VSS.n106 VSS.n80 101.555
R3193 VSS.n566 VSS.n565 97.73
R3194 VSS.n102 VSS.n96 97.5005
R3195 VSS.n1159 VSS.n102 97.5005
R3196 VSS.n1160 VSS.n95 97.5005
R3197 VSS.n1161 VSS.n1160 97.5005
R3198 VSS.n1167 VSS.n1166 97.5005
R3199 VSS.n1168 VSS.n1167 97.5005
R3200 VSS.n650 VSS.n644 97.5005
R3201 VSS.n1148 VSS.n650 97.5005
R3202 VSS.n1149 VSS.n643 97.5005
R3203 VSS.n1150 VSS.n1149 97.5005
R3204 VSS.n1156 VSS.n1155 97.5005
R3205 VSS.n1157 VSS.n1156 97.5005
R3206 VSS.n665 VSS.n659 97.5005
R3207 VSS.n1137 VSS.n665 97.5005
R3208 VSS.n1138 VSS.n658 97.5005
R3209 VSS.n1139 VSS.n1138 97.5005
R3210 VSS.n1145 VSS.n1144 97.5005
R3211 VSS.n1146 VSS.n1145 97.5005
R3212 VSS.n680 VSS.n674 97.5005
R3213 VSS.n1126 VSS.n680 97.5005
R3214 VSS.n1127 VSS.n673 97.5005
R3215 VSS.n1128 VSS.n1127 97.5005
R3216 VSS.n1134 VSS.n1133 97.5005
R3217 VSS.n1135 VSS.n1134 97.5005
R3218 VSS.n695 VSS.n689 97.5005
R3219 VSS.n1115 VSS.n695 97.5005
R3220 VSS.n1116 VSS.n688 97.5005
R3221 VSS.n1117 VSS.n1116 97.5005
R3222 VSS.n1123 VSS.n1122 97.5005
R3223 VSS.n1124 VSS.n1123 97.5005
R3224 VSS.n710 VSS.n704 97.5005
R3225 VSS.n1104 VSS.n710 97.5005
R3226 VSS.n1105 VSS.n703 97.5005
R3227 VSS.n1106 VSS.n1105 97.5005
R3228 VSS.n1112 VSS.n1111 97.5005
R3229 VSS.n1113 VSS.n1112 97.5005
R3230 VSS.n725 VSS.n719 97.5005
R3231 VSS.n1093 VSS.n725 97.5005
R3232 VSS.n1094 VSS.n718 97.5005
R3233 VSS.n1095 VSS.n1094 97.5005
R3234 VSS.n1101 VSS.n1100 97.5005
R3235 VSS.n1102 VSS.n1101 97.5005
R3236 VSS.n786 VSS.n782 97.5005
R3237 VSS.n802 VSS.n786 97.5005
R3238 VSS.n804 VSS.n803 97.5005
R3239 VSS.n805 VSS.n804 97.5005
R3240 VSS.n796 VSS.n795 97.5005
R3241 VSS.n796 VSS.n726 97.5005
R3242 VSS.n833 VSS.n832 96.5764
R3243 VSS.t129 VSS.t319 93.7535
R3244 VSS.t317 VSS.t129 93.7535
R3245 VSS.t339 VSS.t317 93.7535
R3246 VSS.t61 VSS.t138 93.7535
R3247 VSS.t138 VSS.t45 93.7535
R3248 VSS.t45 VSS.t204 93.7535
R3249 VSS.t365 VSS.t179 93.7535
R3250 VSS.n509 VSS.n489 90.2747
R3251 VSS.n862 VSS.t303 86.9189
R3252 VSS.n1065 VSS.t170 86.9189
R3253 VSS.n1031 VSS.t212 86.9189
R3254 VSS.n987 VSS.t207 86.9189
R3255 VSS.n953 VSS.t33 86.9189
R3256 VSS.n909 VSS.t76 86.9189
R3257 VSS.t266 VSS.n108 86.9189
R3258 VSS.n810 VSS.t376 84.5161
R3259 VSS.n788 VSS.t242 84.5161
R3260 VSS.n791 VSS.t119 84.5161
R3261 VSS.n722 VSS.t485 84.5161
R3262 VSS.n714 VSS.t148 84.5161
R3263 VSS.n707 VSS.t412 84.5161
R3264 VSS.n699 VSS.t30 84.5161
R3265 VSS.n692 VSS.t178 84.5161
R3266 VSS.n684 VSS.t117 84.5161
R3267 VSS.n677 VSS.t417 84.5161
R3268 VSS.n669 VSS.t495 84.5161
R3269 VSS.n662 VSS.t224 84.5161
R3270 VSS.n654 VSS.t259 84.5161
R3271 VSS.n647 VSS.t306 84.5161
R3272 VSS.n639 VSS.t196 84.5161
R3273 VSS.n99 VSS.t261 84.5161
R3274 VSS.n303 VSS.t502 84.1574
R3275 VSS.n304 VSS.t96 84.1574
R3276 VSS.n316 VSS.t198 84.1574
R3277 VSS.n317 VSS.t520 84.1574
R3278 VSS.n329 VSS.t540 84.1574
R3279 VSS.n330 VSS.t222 84.1574
R3280 VSS.n342 VSS.t362 84.1574
R3281 VSS.n343 VSS.t327 84.1574
R3282 VSS.n355 VSS.t123 84.1574
R3283 VSS.n356 VSS.t6 84.1574
R3284 VSS.n368 VSS.t44 84.1574
R3285 VSS.n369 VSS.t121 84.1574
R3286 VSS.n381 VSS.t325 84.1574
R3287 VSS.n382 VSS.t518 84.1574
R3288 VSS.n394 VSS.t200 84.1574
R3289 VSS.n395 VSS.t220 84.1574
R3290 VSS.n407 VSS.t230 84.1574
R3291 VSS.n408 VSS.t234 84.1574
R3292 VSS.n420 VSS.t232 84.1574
R3293 VSS.n421 VSS.t228 84.1574
R3294 VSS.n433 VSS.t59 84.1574
R3295 VSS.n434 VSS.t11 84.1574
R3296 VSS.n446 VSS.t184 84.1574
R3297 VSS.n447 VSS.t275 84.1574
R3298 VSS.n459 VSS.t144 84.1574
R3299 VSS.n462 VSS.t314 84.1574
R3300 VSS.n207 VSS.t446 84.1574
R3301 VSS.n200 VSS.t516 84.1574
R3302 VSS.n537 VSS.t425 84.1574
R3303 VSS.n543 VSS.t433 84.1574
R3304 VSS.n545 VSS.t439 84.1574
R3305 VSS.n528 VSS.t17 84.1574
R3306 VSS.n493 VSS.t19 84.1574
R3307 VSS.n496 VSS.t21 84.1574
R3308 VSS.n503 VSS.t23 84.1574
R3309 VSS.n506 VSS.t538 84.1574
R3310 VSS.n836 VSS.t75 83.0558
R3311 VSS.t84 VSS.n862 83.0558
R3312 VSS.t334 VSS.n872 83.0558
R3313 VSS.t237 VSS.n1065 83.0558
R3314 VSS.n1070 VSS.t53 83.0558
R3315 VSS.t359 VSS.n1031 83.0558
R3316 VSS.n1036 VSS.t60 83.0558
R3317 VSS.t551 VSS.n987 83.0558
R3318 VSS.n992 VSS.t488 83.0558
R3319 VSS.t363 VSS.n953 83.0558
R3320 VSS.n958 VSS.t566 83.0558
R3321 VSS.t132 VSS.n909 83.0558
R3322 VSS.n914 VSS.t236 83.0558
R3323 VSS.n108 VSS.t292 83.0558
R3324 VSS.n1171 VSS.t498 83.0558
R3325 VSS.n840 VSS.n741 79.7072
R3326 VSS.n868 VSS.n860 79.7072
R3327 VSS.n1074 VSS.n1057 79.7072
R3328 VSS.n1040 VSS.n1013 79.7072
R3329 VSS.n996 VSS.n979 79.7072
R3330 VSS.n962 VSS.n935 79.7072
R3331 VSS.n918 VSS.n901 79.7072
R3332 VSS.n1175 VSS.n86 79.7072
R3333 VSS.n834 VSS.n745 73.1255
R3334 VSS.n834 VSS.n833 73.1255
R3335 VSS.n864 VSS.n863 73.1255
R3336 VSS.n865 VSS.n864 73.1255
R3337 VSS.n1067 VSS.n1061 73.1255
R3338 VSS.n1067 VSS.n1066 73.1255
R3339 VSS.n1033 VSS.n1017 73.1255
R3340 VSS.n1033 VSS.n1032 73.1255
R3341 VSS.n989 VSS.n983 73.1255
R3342 VSS.n989 VSS.n988 73.1255
R3343 VSS.n955 VSS.n939 73.1255
R3344 VSS.n955 VSS.n954 73.1255
R3345 VSS.n911 VSS.n905 73.1255
R3346 VSS.n911 VSS.n910 73.1255
R3347 VSS.n104 VSS.n103 73.1255
R3348 VSS.n105 VSS.n104 73.1255
R3349 VSS.n839 VSS.n742 69.4405
R3350 VSS.n869 VSS.n854 69.4405
R3351 VSS.n1073 VSS.n1058 69.4405
R3352 VSS.n1039 VSS.n1014 69.4405
R3353 VSS.n995 VSS.n980 69.4405
R3354 VSS.n961 VSS.n936 69.4405
R3355 VSS.n917 VSS.n902 69.4405
R3356 VSS.n1174 VSS.n87 69.4405
R3357 VSS.n301 VSS.n298 68.7561
R3358 VSS.n539 VSS.n536 68.7561
R3359 VSS.n508 VSS.n490 68.7561
R3360 VSS.n569 VSS.n201 68.7561
R3361 VSS.n811 VSS.n783 67.1161
R3362 VSS.n789 VSS.n787 67.1161
R3363 VSS.n792 VSS.n790 67.1161
R3364 VSS.n721 VSS.n720 67.1161
R3365 VSS.n715 VSS.n713 67.1161
R3366 VSS.n706 VSS.n705 67.1161
R3367 VSS.n700 VSS.n698 67.1161
R3368 VSS.n691 VSS.n690 67.1161
R3369 VSS.n685 VSS.n683 67.1161
R3370 VSS.n676 VSS.n675 67.1161
R3371 VSS.n670 VSS.n668 67.1161
R3372 VSS.n661 VSS.n660 67.1161
R3373 VSS.n655 VSS.n653 67.1161
R3374 VSS.n646 VSS.n645 67.1161
R3375 VSS.n640 VSS.n638 67.1161
R3376 VSS.n98 VSS.n97 67.1161
R3377 VSS.n816 VSS.n777 66.9639
R3378 VSS.n817 VSS.n776 66.9639
R3379 VSS.n821 VSS.n818 66.9639
R3380 VSS.n820 VSS.n819 66.9639
R3381 VSS.n771 VSS.n755 66.9639
R3382 VSS.n770 VSS.n756 66.9639
R3383 VSS.n760 VSS.n757 66.9639
R3384 VSS.n759 VSS.n758 66.9639
R3385 VSS.n1242 VSS.n2 66.9639
R3386 VSS.n1241 VSS.n3 66.9639
R3387 VSS.n5 VSS.n4 66.9639
R3388 VSS.n8 VSS.n7 66.9639
R3389 VSS.n19 VSS.n18 66.9639
R3390 VSS.n20 VSS.n17 66.9639
R3391 VSS.n1228 VSS.n21 66.9639
R3392 VSS.n1227 VSS.n22 66.9639
R3393 VSS.n1224 VSS.n24 66.9639
R3394 VSS.n1223 VSS.n25 66.9639
R3395 VSS.n27 VSS.n26 66.9639
R3396 VSS.n30 VSS.n29 66.9639
R3397 VSS.n41 VSS.n40 66.9639
R3398 VSS.n42 VSS.n39 66.9639
R3399 VSS.n1210 VSS.n43 66.9639
R3400 VSS.n1209 VSS.n44 66.9639
R3401 VSS.n1206 VSS.n46 66.9639
R3402 VSS.n1205 VSS.n47 66.9639
R3403 VSS.n49 VSS.n48 66.9639
R3404 VSS.n52 VSS.n51 66.9639
R3405 VSS.n63 VSS.n62 66.9639
R3406 VSS.n64 VSS.n61 66.9639
R3407 VSS.n1192 VSS.n65 66.9639
R3408 VSS.n1191 VSS.n66 66.9639
R3409 VSS.n1188 VSS.n68 66.9639
R3410 VSS.n1187 VSS.n69 66.9639
R3411 VSS.n71 VSS.n70 66.9639
R3412 VSS.n75 VSS.n74 66.9639
R3413 VSS.n117 VSS.n116 66.9639
R3414 VSS.n119 VSS.n118 66.9639
R3415 VSS.n124 VSS.n123 66.9639
R3416 VSS.n125 VSS.n122 66.9639
R3417 VSS.n134 VSS.n133 66.9639
R3418 VSS.n135 VSS.n132 66.9639
R3419 VSS.n613 VSS.n136 66.9639
R3420 VSS.n612 VSS.n137 66.9639
R3421 VSS.n609 VSS.n139 66.9639
R3422 VSS.n608 VSS.n140 66.9639
R3423 VSS.n142 VSS.n141 66.9639
R3424 VSS.n145 VSS.n144 66.9639
R3425 VSS.n160 VSS.n159 66.9639
R3426 VSS.n161 VSS.n158 66.9639
R3427 VSS.n597 VSS.n162 66.9639
R3428 VSS.n596 VSS.n163 66.9639
R3429 VSS.n593 VSS.n165 66.9639
R3430 VSS.n592 VSS.n166 66.9639
R3431 VSS.n168 VSS.n167 66.9639
R3432 VSS.n171 VSS.n170 66.9639
R3433 VSS.n186 VSS.n185 66.9639
R3434 VSS.n187 VSS.n184 66.9639
R3435 VSS.n581 VSS.n188 66.9639
R3436 VSS.n580 VSS.n189 66.9639
R3437 VSS.n577 VSS.n191 66.9639
R3438 VSS.n576 VSS.n192 66.9639
R3439 VSS.n194 VSS.n193 66.9639
R3440 VSS.n198 VSS.n197 66.9639
R3441 VSS.n803 VSS.n785 66.4894
R3442 VSS.n1099 VSS.n718 66.4894
R3443 VSS.n1110 VSS.n703 66.4894
R3444 VSS.n1121 VSS.n688 66.4894
R3445 VSS.n1132 VSS.n673 66.4894
R3446 VSS.n1143 VSS.n658 66.4894
R3447 VSS.n1154 VSS.n643 66.4894
R3448 VSS.n1165 VSS.n95 66.4894
R3449 VSS.n1169 VSS.n92 63.6661
R3450 VSS.t131 VSS.n842 59.8776
R3451 VSS.n866 VSS.t455 59.8776
R3452 VSS.t97 VSS.n1076 59.8776
R3453 VSS.t300 VSS.n1042 59.8776
R3454 VSS.t524 VSS.n998 59.8776
R3455 VSS.t463 VSS.n964 59.8776
R3456 VSS.t65 VSS.n920 59.8776
R3457 VSS.t356 VSS.n1177 59.8776
R3458 VSS.n838 VSS.n837 53.1823
R3459 VSS.n837 VSS.n836 53.1823
R3460 VSS.n871 VSS.n870 53.1823
R3461 VSS.n872 VSS.n871 53.1823
R3462 VSS.n1072 VSS.n1071 53.1823
R3463 VSS.n1071 VSS.n1070 53.1823
R3464 VSS.n1038 VSS.n1037 53.1823
R3465 VSS.n1037 VSS.n1036 53.1823
R3466 VSS.n994 VSS.n993 53.1823
R3467 VSS.n993 VSS.n992 53.1823
R3468 VSS.n960 VSS.n959 53.1823
R3469 VSS.n959 VSS.n958 53.1823
R3470 VSS.n916 VSS.n915 53.1823
R3471 VSS.n915 VSS.n914 53.1823
R3472 VSS.n1173 VSS.n1172 53.1823
R3473 VSS.n1172 VSS.n1171 53.1823
R3474 VSS.n307 VSS.n296 49.4227
R3475 VSS.n292 VSS.n291 49.4227
R3476 VSS.n320 VSS.n289 49.4227
R3477 VSS.n285 VSS.n284 49.4227
R3478 VSS.n333 VSS.n282 49.4227
R3479 VSS.n278 VSS.n277 49.4227
R3480 VSS.n346 VSS.n275 49.4227
R3481 VSS.n271 VSS.n270 49.4227
R3482 VSS.n359 VSS.n268 49.4227
R3483 VSS.n264 VSS.n263 49.4227
R3484 VSS.n372 VSS.n261 49.4227
R3485 VSS.n257 VSS.n256 49.4227
R3486 VSS.n385 VSS.n254 49.4227
R3487 VSS.n250 VSS.n249 49.4227
R3488 VSS.n398 VSS.n247 49.4227
R3489 VSS.n243 VSS.n242 49.4227
R3490 VSS.n411 VSS.n240 49.4227
R3491 VSS.n236 VSS.n235 49.4227
R3492 VSS.n424 VSS.n233 49.4227
R3493 VSS.n229 VSS.n228 49.4227
R3494 VSS.n437 VSS.n226 49.4227
R3495 VSS.n222 VSS.n221 49.4227
R3496 VSS.n450 VSS.n219 49.4227
R3497 VSS.n215 VSS.n214 49.4227
R3498 VSS.n465 VSS.n212 49.4227
R3499 VSS.n460 VSS.n206 49.4227
R3500 VSS.n540 VSS.n534 49.4227
R3501 VSS.n532 VSS.n531 49.4227
R3502 VSS.n549 VSS.n548 49.4227
R3503 VSS.n563 VSS.n562 49.4227
R3504 VSS.n492 VSS.n481 49.4227
R3505 VSS.n499 VSS.n498 49.4227
R3506 VSS.n500 VSS.n491 49.4227
R3507 VSS.n474 VSS.n473 49.4227
R3508 VSS.n841 VSS.n840 48.7505
R3509 VSS.n842 VSS.n841 48.7505
R3510 VSS.n868 VSS.n867 48.7505
R3511 VSS.n867 VSS.n866 48.7505
R3512 VSS.n1075 VSS.n1074 48.7505
R3513 VSS.n1076 VSS.n1075 48.7505
R3514 VSS.n1041 VSS.n1040 48.7505
R3515 VSS.n1042 VSS.n1041 48.7505
R3516 VSS.n997 VSS.n996 48.7505
R3517 VSS.n998 VSS.n997 48.7505
R3518 VSS.n963 VSS.n962 48.7505
R3519 VSS.n964 VSS.n963 48.7505
R3520 VSS.n919 VSS.n918 48.7505
R3521 VSS.n920 VSS.n919 48.7505
R3522 VSS.n1176 VSS.n1175 48.7505
R3523 VSS.n1177 VSS.n1176 48.7505
R3524 VSS.n745 VSS.n741 48.2672
R3525 VSS.n863 VSS.n860 48.2672
R3526 VSS.n1061 VSS.n1057 48.2672
R3527 VSS.n1017 VSS.n1013 48.2672
R3528 VSS.n983 VSS.n979 48.2672
R3529 VSS.n939 VSS.n935 48.2672
R3530 VSS.n905 VSS.n901 48.2672
R3531 VSS.n103 VSS.n86 48.2672
R3532 VSS.n831 VSS.t168 47.9424
R3533 VSS.t179 VSS.n831 45.8116
R3534 VSS.n835 VSS.n743 45.0005
R3535 VSS.n835 VSS.n738 45.0005
R3536 VSS.n859 VSS.n857 45.0005
R3537 VSS.n857 VSS.n856 45.0005
R3538 VSS.n1068 VSS.n1059 45.0005
R3539 VSS.n1068 VSS.n1054 45.0005
R3540 VSS.n1034 VSS.n1015 45.0005
R3541 VSS.n1034 VSS.n1010 45.0005
R3542 VSS.n990 VSS.n981 45.0005
R3543 VSS.n990 VSS.n976 45.0005
R3544 VSS.n956 VSS.n937 45.0005
R3545 VSS.n956 VSS.n932 45.0005
R3546 VSS.n912 VSS.n903 45.0005
R3547 VSS.n912 VSS.n898 45.0005
R3548 VSS.n90 VSS.n88 45.0005
R3549 VSS.n90 VSS.n83 45.0005
R3550 VSS.t537 VSS.n509 43.5008
R3551 VSS.n832 VSS.t365 39.4194
R3552 VSS.n736 VSS.n735 39.0005
R3553 VSS.n828 VSS.n736 39.0005
R3554 VSS.n1088 VSS.n1087 39.0005
R3555 VSS.n1089 VSS.n1088 39.0005
R3556 VSS.n1052 VSS.n875 39.0005
R3557 VSS.n1062 VSS.n1052 39.0005
R3558 VSS.n1008 VSS.n878 39.0005
R3559 VSS.n1028 VSS.n1008 39.0005
R3560 VSS.n974 VSS.n881 39.0005
R3561 VSS.n984 VSS.n974 39.0005
R3562 VSS.n930 VSS.n884 39.0005
R3563 VSS.n950 VSS.n930 39.0005
R3564 VSS.n896 VSS.n887 39.0005
R3565 VSS.n906 VSS.n896 39.0005
R3566 VSS.n81 VSS.n80 39.0005
R3567 VSS.n109 VSS.n81 39.0005
R3568 VSS.n919 VSS.n900 34.4755
R3569 VSS.n963 VSS.n934 34.4755
R3570 VSS.n997 VSS.n978 34.4755
R3571 VSS.n1041 VSS.n1012 34.4755
R3572 VSS.n1075 VSS.n1056 34.4755
R3573 VSS.n867 VSS.n858 34.4755
R3574 VSS.n1176 VSS.n85 34.4755
R3575 VSS.n841 VSS.n740 34.4755
R3576 VSS.n780 VSS.t169 31.7728
R3577 VSS.n850 VSS.t304 31.7728
R3578 VSS.n1082 VSS.t171 31.7728
R3579 VSS.n1048 VSS.t213 31.7728
R3580 VSS.n1004 VSS.t208 31.7728
R3581 VSS.n970 VSS.t34 31.7728
R3582 VSS.n926 VSS.t77 31.7728
R3583 VSS.n892 VSS.t267 31.7728
R3584 VSS.n615 VSS.n130 28.8579
R3585 VSS.n606 VSS.n143 28.8579
R3586 VSS.n599 VSS.n156 28.8579
R3587 VSS.n590 VSS.n169 28.8579
R3588 VSS.n583 VSS.n182 28.8579
R3589 VSS.n574 VSS.n195 28.8579
R3590 VSS.n1194 VSS.n59 28.8579
R3591 VSS.n1203 VSS.n50 28.8579
R3592 VSS.n1212 VSS.n37 28.8579
R3593 VSS.n1221 VSS.n28 28.8579
R3594 VSS.n1230 VSS.n15 28.8579
R3595 VSS.n1239 VSS.n6 28.8579
R3596 VSS.n768 VSS.n761 28.8579
R3597 VSS.n823 VSS.n774 28.8579
R3598 VSS.n1185 VSS.n72 28.8579
R3599 VSS.n622 VSS.n121 28.857
R3600 VSS.n127 VSS.n121 28.6936
R3601 VSS.n629 VSS.n72 28.6927
R3602 VSS.n516 VSS.n195 28.6927
R3603 VSS.n510 VSS.n182 28.6927
R3604 VSS.n179 VSS.n169 28.6927
R3605 VSS.n174 VSS.n156 28.6927
R3606 VSS.n153 VSS.n143 28.6927
R3607 VSS.n148 VSS.n130 28.6927
R3608 VSS.n800 VSS.n774 28.6927
R3609 VSS.n747 VSS.n6 28.6927
R3610 VSS.n1021 VSS.n28 28.6927
R3611 VSS.n943 VSS.n50 28.6927
R3612 VSS.n110 VSS.n59 28.6927
R3613 VSS.n940 VSS.n37 28.6927
R3614 VSS.n1018 VSS.n15 28.6927
R3615 VSS.n764 VSS.n761 28.6927
R3616 VSS.n779 VSS.n778 25.9728
R3617 VSS.n734 VSS.n733 25.9728
R3618 VSS.n851 VSS.n849 25.9728
R3619 VSS.n852 VSS.n848 25.9728
R3620 VSS.n1081 VSS.n876 25.9728
R3621 VSS.n1080 VSS.n877 25.9728
R3622 VSS.n1047 VSS.n879 25.9728
R3623 VSS.n1046 VSS.n880 25.9728
R3624 VSS.n1003 VSS.n882 25.9728
R3625 VSS.n1002 VSS.n883 25.9728
R3626 VSS.n969 VSS.n885 25.9728
R3627 VSS.n968 VSS.n886 25.9728
R3628 VSS.n925 VSS.n888 25.9728
R3629 VSS.n924 VSS.n889 25.9728
R3630 VSS.n891 VSS.n890 25.9728
R3631 VSS.n79 VSS.n78 25.9728
R3632 VSS.n842 VSS.n738 23.1787
R3633 VSS.n866 VSS.n856 23.1787
R3634 VSS.n1076 VSS.n1054 23.1787
R3635 VSS.n1042 VSS.n1010 23.1787
R3636 VSS.n998 VSS.n976 23.1787
R3637 VSS.n964 VSS.n932 23.1787
R3638 VSS.n920 VSS.n898 23.1787
R3639 VSS.n1177 VSS.n83 23.1787
R3640 VSS.n829 VSS.n741 23.1494
R3641 VSS.n860 VSS.n731 23.1494
R3642 VSS.n1063 VSS.n1057 23.1494
R3643 VSS.n1029 VSS.n1013 23.1494
R3644 VSS.n985 VSS.n979 23.1494
R3645 VSS.n951 VSS.n935 23.1494
R3646 VSS.n907 VSS.n901 23.1494
R3647 VSS.n106 VSS.n86 23.1494
R3648 VSS.n82 VSS.n77 22.5005
R3649 VSS.n91 VSS.n82 22.5005
R3650 VSS.n737 VSS.n732 22.5005
R3651 VSS.n737 VSS.n727 22.5005
R3652 VSS.n1085 VSS.n874 22.5005
R3653 VSS.n874 VSS.n873 22.5005
R3654 VSS.n1053 VSS.n1051 22.5005
R3655 VSS.n1069 VSS.n1053 22.5005
R3656 VSS.n1009 VSS.n1007 22.5005
R3657 VSS.n1035 VSS.n1009 22.5005
R3658 VSS.n975 VSS.n973 22.5005
R3659 VSS.n991 VSS.n975 22.5005
R3660 VSS.n931 VSS.n929 22.5005
R3661 VSS.n957 VSS.n931 22.5005
R3662 VSS.n897 VSS.n895 22.5005
R3663 VSS.n913 VSS.n897 22.5005
R3664 VSS.n1162 VSS.n1161 19.761
R3665 VSS.n1151 VSS.n1150 19.761
R3666 VSS.n1140 VSS.n1139 19.761
R3667 VSS.n1129 VSS.n1128 19.761
R3668 VSS.n1118 VSS.n1117 19.761
R3669 VSS.n1107 VSS.n1106 19.761
R3670 VSS.n1096 VSS.n1095 19.761
R3671 VSS.n806 VSS.n805 19.761
R3672 VSS.n1170 VSS.n91 19.4911
R3673 VSS.n540 VSS.n539 19.3338
R3674 VSS.n541 VSS.n540 19.3338
R3675 VSS.n541 VSS.n531 19.3338
R3676 VSS.n547 VSS.n531 19.3338
R3677 VSS.n548 VSS.n547 19.3338
R3678 VSS.n548 VSS.n479 19.3338
R3679 VSS.n562 VSS.n479 19.3338
R3680 VSS.n562 VSS.n561 19.3338
R3681 VSS.n561 VSS.n481 19.3338
R3682 VSS.n484 VSS.n481 19.3338
R3683 VSS.n499 VSS.n484 19.3338
R3684 VSS.n501 VSS.n499 19.3338
R3685 VSS.n501 VSS.n500 19.3338
R3686 VSS.n500 VSS.n490 19.3338
R3687 VSS.n301 VSS.n296 19.3338
R3688 VSS.n296 VSS.n295 19.3338
R3689 VSS.n295 VSS.n291 19.3338
R3690 VSS.n314 VSS.n291 19.3338
R3691 VSS.n314 VSS.n289 19.3338
R3692 VSS.n289 VSS.n288 19.3338
R3693 VSS.n288 VSS.n284 19.3338
R3694 VSS.n327 VSS.n284 19.3338
R3695 VSS.n327 VSS.n282 19.3338
R3696 VSS.n282 VSS.n281 19.3338
R3697 VSS.n281 VSS.n277 19.3338
R3698 VSS.n340 VSS.n277 19.3338
R3699 VSS.n340 VSS.n275 19.3338
R3700 VSS.n275 VSS.n274 19.3338
R3701 VSS.n274 VSS.n270 19.3338
R3702 VSS.n353 VSS.n270 19.3338
R3703 VSS.n353 VSS.n268 19.3338
R3704 VSS.n268 VSS.n267 19.3338
R3705 VSS.n267 VSS.n263 19.3338
R3706 VSS.n366 VSS.n263 19.3338
R3707 VSS.n366 VSS.n261 19.3338
R3708 VSS.n261 VSS.n260 19.3338
R3709 VSS.n260 VSS.n256 19.3338
R3710 VSS.n379 VSS.n256 19.3338
R3711 VSS.n379 VSS.n254 19.3338
R3712 VSS.n254 VSS.n253 19.3338
R3713 VSS.n253 VSS.n249 19.3338
R3714 VSS.n392 VSS.n249 19.3338
R3715 VSS.n392 VSS.n247 19.3338
R3716 VSS.n247 VSS.n246 19.3338
R3717 VSS.n246 VSS.n242 19.3338
R3718 VSS.n405 VSS.n242 19.3338
R3719 VSS.n405 VSS.n240 19.3338
R3720 VSS.n240 VSS.n239 19.3338
R3721 VSS.n239 VSS.n235 19.3338
R3722 VSS.n418 VSS.n235 19.3338
R3723 VSS.n418 VSS.n233 19.3338
R3724 VSS.n233 VSS.n232 19.3338
R3725 VSS.n232 VSS.n228 19.3338
R3726 VSS.n431 VSS.n228 19.3338
R3727 VSS.n431 VSS.n226 19.3338
R3728 VSS.n226 VSS.n225 19.3338
R3729 VSS.n225 VSS.n221 19.3338
R3730 VSS.n444 VSS.n221 19.3338
R3731 VSS.n444 VSS.n219 19.3338
R3732 VSS.n219 VSS.n218 19.3338
R3733 VSS.n218 VSS.n214 19.3338
R3734 VSS.n457 VSS.n214 19.3338
R3735 VSS.n457 VSS.n212 19.3338
R3736 VSS.n212 VSS.n211 19.3338
R3737 VSS.n211 VSS.n206 19.3338
R3738 VSS.n472 VSS.n206 19.3338
R3739 VSS.n473 VSS.n472 19.3338
R3740 VSS.n473 VSS.n201 19.3338
R3741 VSS.n742 VSS.n732 18.2672
R3742 VSS.n1085 VSS.n854 18.2672
R3743 VSS.n1058 VSS.n1051 18.2672
R3744 VSS.n1014 VSS.n1007 18.2672
R3745 VSS.n980 VSS.n973 18.2672
R3746 VSS.n936 VSS.n929 18.2672
R3747 VSS.n902 VSS.n895 18.2672
R3748 VSS.n87 VSS.n77 18.2672
R3749 VSS.n777 VSS.t320 17.4005
R3750 VSS.n777 VSS.t130 17.4005
R3751 VSS.n776 VSS.t318 17.4005
R3752 VSS.n776 VSS.t340 17.4005
R3753 VSS.n818 VSS.t62 17.4005
R3754 VSS.n818 VSS.t139 17.4005
R3755 VSS.n819 VSS.t46 17.4005
R3756 VSS.n819 VSS.t205 17.4005
R3757 VSS.n755 VSS.t312 17.4005
R3758 VSS.n755 VSS.t454 17.4005
R3759 VSS.n756 VSS.t457 17.4005
R3760 VSS.n756 VSS.t251 17.4005
R3761 VSS.n757 VSS.t336 17.4005
R3762 VSS.n757 VSS.t128 17.4005
R3763 VSS.n758 VSS.t269 17.4005
R3764 VSS.n758 VSS.t368 17.4005
R3765 VSS.n2 VSS.t99 17.4005
R3766 VSS.n2 VSS.t52 17.4005
R3767 VSS.n3 VSS.t404 17.4005
R3768 VSS.n3 VSS.t69 17.4005
R3769 VSS.n4 VSS.t331 17.4005
R3770 VSS.n4 VSS.t542 17.4005
R3771 VSS.n7 VSS.t329 17.4005
R3772 VSS.n7 VSS.t544 17.4005
R3773 VSS.n18 VSS.t490 17.4005
R3774 VSS.n18 VSS.t298 17.4005
R3775 VSS.n17 VSS.t150 17.4005
R3776 VSS.n17 VSS.t374 17.4005
R3777 VSS.n21 VSS.t83 17.4005
R3778 VSS.n21 VSS.t80 17.4005
R3779 VSS.n22 VSS.t146 17.4005
R3780 VSS.n22 VSS.t295 17.4005
R3781 VSS.n24 VSS.t512 17.4005
R3782 VSS.n24 VSS.t396 17.4005
R3783 VSS.n25 VSS.t394 17.4005
R3784 VSS.n25 VSS.t398 17.4005
R3785 VSS.n26 VSS.t289 17.4005
R3786 VSS.n26 VSS.t574 17.4005
R3787 VSS.n29 VSS.t577 17.4005
R3788 VSS.n29 VSS.t431 17.4005
R3789 VSS.n40 VSS.t461 17.4005
R3790 VSS.n40 VSS.t467 17.4005
R3791 VSS.n39 VSS.t459 17.4005
R3792 VSS.n39 VSS.t465 17.4005
R3793 VSS.n43 VSS.t410 17.4005
R3794 VSS.n43 VSS.t568 17.4005
R3795 VSS.n44 VSS.t408 17.4005
R3796 VSS.n44 VSS.t392 17.4005
R3797 VSS.n46 VSS.t64 17.4005
R3798 VSS.n46 VSS.t88 17.4005
R3799 VSS.n47 VSS.t570 17.4005
R3800 VSS.n47 VSS.t557 17.4005
R3801 VSS.n48 VSS.t254 17.4005
R3802 VSS.n48 VSS.t182 17.4005
R3803 VSS.n51 VSS.t422 17.4005
R3804 VSS.n51 VSS.t71 17.4005
R3805 VSS.n62 VSS.t190 17.4005
R3806 VSS.n62 VSS.t526 17.4005
R3807 VSS.n61 VSS.t160 17.4005
R3808 VSS.n61 VSS.t497 17.4005
R3809 VSS.n65 VSS.t355 17.4005
R3810 VSS.n65 VSS.t492 17.4005
R3811 VSS.n66 VSS.t487 17.4005
R3812 VSS.n66 VSS.t283 17.4005
R3813 VSS.n68 VSS.t240 17.4005
R3814 VSS.n68 VSS.t265 17.4005
R3815 VSS.n69 VSS.t218 17.4005
R3816 VSS.n69 VSS.t561 17.4005
R3817 VSS.n70 VSS.t479 17.4005
R3818 VSS.n70 VSS.t273 17.4005
R3819 VSS.n74 VSS.t104 17.4005
R3820 VSS.n74 VSS.t257 17.4005
R3821 VSS.n116 VSS.t156 17.4005
R3822 VSS.n116 VSS.t444 17.4005
R3823 VSS.n118 VSS.t158 17.4005
R3824 VSS.n118 VSS.t167 17.4005
R3825 VSS.n123 VSS.t427 17.4005
R3826 VSS.n123 VSS.t475 17.4005
R3827 VSS.n122 VSS.t192 17.4005
R3828 VSS.n122 VSS.t535 17.4005
R3829 VSS.n133 VSS.t370 17.4005
R3830 VSS.n133 VSS.t25 17.4005
R3831 VSS.n132 VSS.t506 17.4005
R3832 VSS.n132 VSS.t215 17.4005
R3833 VSS.n136 VSS.t115 17.4005
R3834 VSS.n136 VSS.t350 17.4005
R3835 VSS.n137 VSS.t437 17.4005
R3836 VSS.n137 VSS.t435 17.4005
R3837 VSS.n139 VSS.t406 17.4005
R3838 VSS.n139 VSS.t548 17.4005
R3839 VSS.n140 VSS.t550 17.4005
R3840 VSS.n140 VSS.t55 17.4005
R3841 VSS.n141 VSS.t533 17.4005
R3842 VSS.n141 VSS.t287 17.4005
R3843 VSS.n144 VSS.t400 17.4005
R3844 VSS.n144 VSS.t101 17.4005
R3845 VSS.n159 VSS.t358 17.4005
R3846 VSS.n159 VSS.t448 17.4005
R3847 VSS.n158 VSS.t285 17.4005
R3848 VSS.n158 VSS.t106 17.4005
R3849 VSS.n162 VSS.t402 17.4005
R3850 VSS.n162 VSS.t450 17.4005
R3851 VSS.n163 VSS.t528 17.4005
R3852 VSS.n163 VSS.t137 17.4005
R3853 VSS.n165 VSS.t154 17.4005
R3854 VSS.n165 VSS.t563 17.4005
R3855 VSS.n166 VSS.t583 17.4005
R3856 VSS.n166 VSS.t580 17.4005
R3857 VSS.n167 VSS.t514 17.4005
R3858 VSS.n167 VSS.t508 17.4005
R3859 VSS.n170 VSS.t429 17.4005
R3860 VSS.n170 VSS.t316 17.4005
R3861 VSS.n185 VSS.t141 17.4005
R3862 VSS.n185 VSS.t176 17.4005
R3863 VSS.n184 VSS.t94 17.4005
R3864 VSS.n184 VSS.t49 17.4005
R3865 VSS.n188 VSS.t477 17.4005
R3866 VSS.n188 VSS.t291 17.4005
R3867 VSS.n189 VSS.t67 17.4005
R3868 VSS.n189 VSS.t92 17.4005
R3869 VSS.n191 VSS.t572 17.4005
R3870 VSS.n191 VSS.t40 17.4005
R3871 VSS.n192 VSS.t310 17.4005
R3872 VSS.n192 VSS.t452 17.4005
R3873 VSS.n193 VSS.t194 17.4005
R3874 VSS.n193 VSS.t500 17.4005
R3875 VSS.n197 VSS.t323 17.4005
R3876 VSS.n197 VSS.t90 17.4005
R3877 VSS.n783 VSS.t379 17.4005
R3878 VSS.n783 VSS.t565 17.4005
R3879 VSS.n787 VSS.t226 17.4005
R3880 VSS.n787 VSS.t442 17.4005
R3881 VSS.n790 VSS.t388 17.4005
R3882 VSS.n790 VSS.t15 17.4005
R3883 VSS.n720 VSS.t390 17.4005
R3884 VSS.n720 VSS.t384 17.4005
R3885 VSS.n713 VSS.t113 17.4005
R3886 VSS.n713 VSS.t510 17.4005
R3887 VSS.n705 VSS.t125 17.4005
R3888 VSS.n705 VSS.t346 17.4005
R3889 VSS.n698 VSS.t471 17.4005
R3890 VSS.n698 VSS.t554 17.4005
R3891 VSS.n690 VSS.t483 17.4005
R3892 VSS.n690 VSS.t473 17.4005
R3893 VSS.n683 VSS.t1 17.4005
R3894 VSS.n683 VSS.t244 17.4005
R3895 VSS.n675 VSS.t271 17.4005
R3896 VSS.n675 VSS.t165 17.4005
R3897 VSS.n668 VSS.t420 17.4005
R3898 VSS.n668 VSS.t279 17.4005
R3899 VSS.n660 VSS.t173 17.4005
R3900 VSS.n660 VSS.t530 17.4005
R3901 VSS.n653 VSS.t344 17.4005
R3902 VSS.n653 VSS.t559 17.4005
R3903 VSS.n645 VSS.t8 17.4005
R3904 VSS.n645 VSS.t152 17.4005
R3905 VSS.n638 VSS.t263 17.4005
R3906 VSS.n638 VSS.t210 17.4005
R3907 VSS.n97 VSS.t281 17.4005
R3908 VSS.n97 VSS.t372 17.4005
R3909 VSS.n1164 VSS.n1163 17.2064
R3910 VSS.n1163 VSS.n1162 17.2064
R3911 VSS.n1153 VSS.n1152 17.2064
R3912 VSS.n1152 VSS.n1151 17.2064
R3913 VSS.n1142 VSS.n1141 17.2064
R3914 VSS.n1141 VSS.n1140 17.2064
R3915 VSS.n1131 VSS.n1130 17.2064
R3916 VSS.n1130 VSS.n1129 17.2064
R3917 VSS.n1120 VSS.n1119 17.2064
R3918 VSS.n1119 VSS.n1118 17.2064
R3919 VSS.n1109 VSS.n1108 17.2064
R3920 VSS.n1108 VSS.n1107 17.2064
R3921 VSS.n1098 VSS.n1097 17.2064
R3922 VSS.n1097 VSS.n1096 17.2064
R3923 VSS.n808 VSS.n807 17.2064
R3924 VSS.n807 VSS.n806 17.2064
R3925 VSS.n844 VSS.n843 15.3952
R3926 VSS.n843 VSS.t377 15.3952
R3927 VSS.n1086 VSS.n730 15.3952
R3928 VSS.t216 VSS.n730 15.3952
R3929 VSS.n1078 VSS.n1077 15.3952
R3930 VSS.n1077 VSS.t174 15.3952
R3931 VSS.n1044 VSS.n1043 15.3952
R3932 VSS.n1043 VSS.t78 15.3952
R3933 VSS.n1000 VSS.n999 15.3952
R3934 VSS.n999 VSS.t2 15.3952
R3935 VSS.n966 VSS.n965 15.3952
R3936 VSS.n965 VSS.t255 15.3952
R3937 VSS.n922 VSS.n921 15.3952
R3938 VSS.n921 VSS.t110 15.3952
R3939 VSS.n1179 VSS.n1178 15.3952
R3940 VSS.n1178 VSS.t308 15.3952
R3941 VSS.n801 VSS.n800 12.785
R3942 VSS.n828 VSS.n827 10.6543
R3943 VSS.n812 VSS.n782 7.71988
R3944 VSS.n803 VSS.n784 7.71988
R3945 VSS.n795 VSS.n794 7.71988
R3946 VSS.n793 VSS.n719 7.71988
R3947 VSS.n723 VSS.n718 7.71988
R3948 VSS.n1100 VSS.n717 7.71988
R3949 VSS.n716 VSS.n704 7.71988
R3950 VSS.n708 VSS.n703 7.71988
R3951 VSS.n1111 VSS.n702 7.71988
R3952 VSS.n701 VSS.n689 7.71988
R3953 VSS.n693 VSS.n688 7.71988
R3954 VSS.n1122 VSS.n687 7.71988
R3955 VSS.n686 VSS.n674 7.71988
R3956 VSS.n678 VSS.n673 7.71988
R3957 VSS.n1133 VSS.n672 7.71988
R3958 VSS.n671 VSS.n659 7.71988
R3959 VSS.n663 VSS.n658 7.71988
R3960 VSS.n1144 VSS.n657 7.71988
R3961 VSS.n656 VSS.n644 7.71988
R3962 VSS.n648 VSS.n643 7.71988
R3963 VSS.n1155 VSS.n642 7.71988
R3964 VSS.n641 VSS.n96 7.71988
R3965 VSS.n100 VSS.n95 7.71988
R3966 VSS.n1166 VSS.n94 7.71988
R3967 VSS.n297 VSS.n76 5.90952
R3968 VSS.n778 VSS.t180 5.8005
R3969 VSS.n778 VSS.t366 5.8005
R3970 VSS.n733 VSS.t414 5.8005
R3971 VSS.n733 VSS.t36 5.8005
R3972 VSS.n849 VSS.t85 5.8005
R3973 VSS.n849 VSS.t32 5.8005
R3974 VSS.n848 VSS.t13 5.8005
R3975 VSS.n848 VSS.t504 5.8005
R3976 VSS.n876 VSS.t238 5.8005
R3977 VSS.n876 VSS.t203 5.8005
R3978 VSS.n877 VSS.t135 5.8005
R3979 VSS.n877 VSS.t481 5.8005
R3980 VSS.n879 VSS.t360 5.8005
R3981 VSS.n879 VSS.t188 5.8005
R3982 VSS.n880 VSS.t302 5.8005
R3983 VSS.n880 VSS.t246 5.8005
R3984 VSS.n882 VSS.t552 5.8005
R3985 VSS.n882 VSS.t38 5.8005
R3986 VSS.n883 VSS.t186 5.8005
R3987 VSS.n883 VSS.t248 5.8005
R3988 VSS.n885 VSS.t364 5.8005
R3989 VSS.n885 VSS.t546 5.8005
R3990 VSS.n886 VSS.t348 5.8005
R3991 VSS.n886 VSS.t277 5.8005
R3992 VSS.n888 VSS.t133 5.8005
R3993 VSS.n888 VSS.t333 5.8005
R3994 VSS.n889 VSS.t74 5.8005
R3995 VSS.n889 VSS.t342 5.8005
R3996 VSS.n890 VSS.t293 5.8005
R3997 VSS.n890 VSS.t353 5.8005
R3998 VSS.n78 VSS.t338 5.8005
R3999 VSS.n78 VSS.t57 5.8005
R4000 VSS.n807 VSS.n797 5.79462
R4001 VSS.n1097 VSS.n712 5.79462
R4002 VSS.n1108 VSS.n697 5.79462
R4003 VSS.n1119 VSS.n682 5.79462
R4004 VSS.n1130 VSS.n667 5.79462
R4005 VSS.n1141 VSS.n652 5.79462
R4006 VSS.n1152 VSS.n637 5.79462
R4007 VSS.n1163 VSS.n93 5.79462
R4008 VSS.n813 VSS.n812 3.89165
R4009 VSS.n836 VSS.n738 3.86354
R4010 VSS.n872 VSS.n856 3.86354
R4011 VSS.n1070 VSS.n1054 3.86354
R4012 VSS.n1036 VSS.n1010 3.86354
R4013 VSS.n992 VSS.n976 3.86354
R4014 VSS.n958 VSS.n932 3.86354
R4015 VSS.n914 VSS.n898 3.86354
R4016 VSS.n1171 VSS.n83 3.86354
R4017 VSS.n1182 VSS.n76 3.78262
R4018 VSS.n571 VSS 3.50128
R4019 VSS.n298 VSS.n297 3.46248
R4020 VSS.n307 VSS.n306 3.46248
R4021 VSS.n292 VSS.n290 3.46248
R4022 VSS.n320 VSS.n319 3.46248
R4023 VSS.n285 VSS.n283 3.46248
R4024 VSS.n333 VSS.n332 3.46248
R4025 VSS.n278 VSS.n276 3.46248
R4026 VSS.n346 VSS.n345 3.46248
R4027 VSS.n271 VSS.n269 3.46248
R4028 VSS.n359 VSS.n358 3.46248
R4029 VSS.n264 VSS.n262 3.46248
R4030 VSS.n372 VSS.n371 3.46248
R4031 VSS.n257 VSS.n255 3.46248
R4032 VSS.n385 VSS.n384 3.46248
R4033 VSS.n250 VSS.n248 3.46248
R4034 VSS.n398 VSS.n397 3.46248
R4035 VSS.n243 VSS.n241 3.46248
R4036 VSS.n411 VSS.n410 3.46248
R4037 VSS.n236 VSS.n234 3.46248
R4038 VSS.n424 VSS.n423 3.46248
R4039 VSS.n229 VSS.n227 3.46248
R4040 VSS.n437 VSS.n436 3.46248
R4041 VSS.n222 VSS.n220 3.46248
R4042 VSS.n450 VSS.n449 3.46248
R4043 VSS.n215 VSS.n213 3.46248
R4044 VSS.n465 VSS.n464 3.46248
R4045 VSS.n461 VSS.n460 3.46248
R4046 VSS.n474 VSS.n205 3.46248
R4047 VSS.n536 VSS.n199 3.46248
R4048 VSS.n534 VSS.n533 3.46248
R4049 VSS.n544 VSS.n532 3.46248
R4050 VSS.n549 VSS.n530 3.46248
R4051 VSS.n563 VSS.n478 3.46248
R4052 VSS.n494 VSS.n492 3.46248
R4053 VSS.n498 VSS.n497 3.46248
R4054 VSS.n504 VSS.n491 3.46248
R4055 VSS.n508 VSS.n507 3.46248
R4056 VSS.n570 VSS.n569 3.46248
R4057 VSS.n623 VSS.n117 3.0154
R4058 VSS VSS.n1182 2.89807
R4059 VSS.n584 VSS.n181 2.768
R4060 VSS.n579 VSS.n183 2.768
R4061 VSS.n594 VSS.n164 2.768
R4062 VSS.n589 VSS.n172 2.768
R4063 VSS.n600 VSS.n155 2.768
R4064 VSS.n595 VSS.n157 2.768
R4065 VSS.n610 VSS.n138 2.768
R4066 VSS.n605 VSS.n146 2.768
R4067 VSS.n616 VSS.n129 2.768
R4068 VSS.n611 VSS.n131 2.768
R4069 VSS.n621 VSS.n126 2.768
R4070 VSS.n578 VSS.n190 2.768
R4071 VSS.n573 VSS.n572 2.768
R4072 VSS.n815 VSS.n775 2.768
R4073 VSS.n824 VSS.n773 2.768
R4074 VSS.n1238 VSS.n9 2.768
R4075 VSS.n1243 VSS.n1 2.768
R4076 VSS.n1220 VSS.n31 2.768
R4077 VSS.n1225 VSS.n23 2.768
R4078 VSS.n1202 VSS.n53 2.768
R4079 VSS.n1207 VSS.n45 2.768
R4080 VSS.n1195 VSS.n58 2.768
R4081 VSS.n1190 VSS.n60 2.768
R4082 VSS.n1213 VSS.n36 2.768
R4083 VSS.n1208 VSS.n38 2.768
R4084 VSS.n1231 VSS.n14 2.768
R4085 VSS.n1226 VSS.n16 2.768
R4086 VSS.n772 VSS.n754 2.768
R4087 VSS.n767 VSS.n0 2.768
R4088 VSS.n1189 VSS.n67 2.768
R4089 VSS.n1184 VSS.n1183 2.768
R4090 VSS.n130 VSS.n128 2.52995
R4091 VSS.n147 VSS.n143 2.52995
R4092 VSS.n156 VSS.n154 2.52995
R4093 VSS.n173 VSS.n169 2.52995
R4094 VSS.n182 VSS.n180 2.52995
R4095 VSS.n513 VSS.n195 2.52995
R4096 VSS.n59 VSS.n57 2.52995
R4097 VSS.n54 VSS.n50 2.52995
R4098 VSS.n37 VSS.n35 2.52995
R4099 VSS.n32 VSS.n28 2.52995
R4100 VSS.n15 VSS.n13 2.52995
R4101 VSS.n10 VSS.n6 2.52995
R4102 VSS.n763 VSS.n761 2.52995
R4103 VSS.n774 VSS.n753 2.52995
R4104 VSS.n630 VSS.n72 2.52995
R4105 VSS.n121 VSS.n115 2.52995
R4106 VSS.n1182 VSS 2.40675
R4107 VSS.n814 VSS.n813 2.3961
R4108 VSS.n539 VSS.n538 2.3255
R4109 VSS.n542 VSS.n541 2.3255
R4110 VSS.n547 VSS.n546 2.3255
R4111 VSS.n529 VSS.n479 2.3255
R4112 VSS.n561 VSS.n480 2.3255
R4113 VSS.n495 VSS.n484 2.3255
R4114 VSS.n502 VSS.n501 2.3255
R4115 VSS.n505 VSS.n490 2.3255
R4116 VSS.n302 VSS.n301 2.3255
R4117 VSS.n305 VSS.n295 2.3255
R4118 VSS.n315 VSS.n314 2.3255
R4119 VSS.n318 VSS.n288 2.3255
R4120 VSS.n328 VSS.n327 2.3255
R4121 VSS.n331 VSS.n281 2.3255
R4122 VSS.n341 VSS.n340 2.3255
R4123 VSS.n344 VSS.n274 2.3255
R4124 VSS.n354 VSS.n353 2.3255
R4125 VSS.n357 VSS.n267 2.3255
R4126 VSS.n367 VSS.n366 2.3255
R4127 VSS.n370 VSS.n260 2.3255
R4128 VSS.n380 VSS.n379 2.3255
R4129 VSS.n383 VSS.n253 2.3255
R4130 VSS.n393 VSS.n392 2.3255
R4131 VSS.n396 VSS.n246 2.3255
R4132 VSS.n406 VSS.n405 2.3255
R4133 VSS.n409 VSS.n239 2.3255
R4134 VSS.n419 VSS.n418 2.3255
R4135 VSS.n422 VSS.n232 2.3255
R4136 VSS.n432 VSS.n431 2.3255
R4137 VSS.n435 VSS.n225 2.3255
R4138 VSS.n445 VSS.n444 2.3255
R4139 VSS.n448 VSS.n218 2.3255
R4140 VSS.n458 VSS.n457 2.3255
R4141 VSS.n463 VSS.n211 2.3255
R4142 VSS.n472 VSS.n208 2.3255
R4143 VSS.n204 VSS.n201 2.3255
R4144 VSS.n813 VSS.n781 2.28621
R4145 VSS.n840 VSS.n839 2.2405
R4146 VSS.n869 VSS.n868 2.2405
R4147 VSS.n1074 VSS.n1073 2.2405
R4148 VSS.n1040 VSS.n1039 2.2405
R4149 VSS.n996 VSS.n995 2.2405
R4150 VSS.n962 VSS.n961 2.2405
R4151 VSS.n918 VSS.n917 2.2405
R4152 VSS.n1175 VSS.n1174 2.2405
R4153 VSS.n833 VSS.t413 1.93202
R4154 VSS.t12 VSS.n865 1.93202
R4155 VSS.n1066 VSS.t134 1.93202
R4156 VSS.n1032 VSS.t301 1.93202
R4157 VSS.n988 VSS.t185 1.93202
R4158 VSS.n954 VSS.t347 1.93202
R4159 VSS.n910 VSS.t73 1.93202
R4160 VSS.n105 VSS.t337 1.93202
R4161 VSS.n846 VSS.n732 1.56378
R4162 VSS.n1085 VSS.n1084 1.56378
R4163 VSS.n1051 VSS.n1050 1.56378
R4164 VSS.n1007 VSS.n1006 1.56378
R4165 VSS.n973 VSS.n972 1.56378
R4166 VSS.n929 VSS.n928 1.56378
R4167 VSS.n895 VSS.n894 1.56378
R4168 VSS.n1181 VSS.n77 1.56378
R4169 VSS VSS.n772 1.3768
R4170 VSS VSS.n1243 1.3768
R4171 VSS.n14 VSS 1.3768
R4172 VSS VSS.n1225 1.3768
R4173 VSS.n36 VSS 1.3768
R4174 VSS VSS.n1207 1.3768
R4175 VSS.n58 VSS 1.3768
R4176 VSS VSS.n1189 1.3768
R4177 VSS.n781 VSS.n735 1.37182
R4178 VSS.n1087 VSS.n847 1.37182
R4179 VSS.n1083 VSS.n875 1.37182
R4180 VSS.n1049 VSS.n878 1.37182
R4181 VSS.n1005 VSS.n881 1.37182
R4182 VSS.n971 VSS.n884 1.37182
R4183 VSS.n927 VSS.n887 1.37182
R4184 VSS.n893 VSS.n80 1.37182
R4185 VSS.n814 VSS 1.17495
R4186 VSS.n846 VSS.n845 0.785098
R4187 VSS.n1084 VSS.n853 0.785098
R4188 VSS.n1079 VSS.n1050 0.785098
R4189 VSS.n1045 VSS.n1006 0.785098
R4190 VSS.n1001 VSS.n972 0.785098
R4191 VSS.n967 VSS.n928 0.785098
R4192 VSS.n923 VSS.n894 0.785098
R4193 VSS.n1181 VSS.n1180 0.785098
R4194 VSS VSS.n793 0.669618
R4195 VSS VSS.n716 0.669618
R4196 VSS VSS.n701 0.669618
R4197 VSS VSS.n686 0.669618
R4198 VSS VSS.n671 0.669618
R4199 VSS VSS.n656 0.669618
R4200 VSS VSS.n641 0.669618
R4201 VSS.n622 VSS.n120 0.58175
R4202 VSS.n615 VSS.n614 0.58175
R4203 VSS.n607 VSS.n606 0.58175
R4204 VSS.n599 VSS.n598 0.58175
R4205 VSS.n591 VSS.n590 0.58175
R4206 VSS.n583 VSS.n582 0.58175
R4207 VSS.n575 VSS.n574 0.58175
R4208 VSS.n809 VSS.n808 0.58175
R4209 VSS.n1098 VSS.n724 0.58175
R4210 VSS.n1109 VSS.n709 0.58175
R4211 VSS.n1120 VSS.n694 0.58175
R4212 VSS.n1131 VSS.n679 0.58175
R4213 VSS.n1142 VSS.n664 0.58175
R4214 VSS.n1153 VSS.n649 0.58175
R4215 VSS.n1164 VSS.n101 0.58175
R4216 VSS.n823 VSS.n822 0.58175
R4217 VSS.n769 VSS.n768 0.58175
R4218 VSS.n1240 VSS.n1239 0.58175
R4219 VSS.n1230 VSS.n1229 0.58175
R4220 VSS.n1222 VSS.n1221 0.58175
R4221 VSS.n1212 VSS.n1211 0.58175
R4222 VSS.n1204 VSS.n1203 0.58175
R4223 VSS.n1194 VSS.n1193 0.58175
R4224 VSS.n1186 VSS.n1185 0.58175
R4225 VSS.n815 VSS.n814 0.53826
R4226 VSS VSS.n846 0.522821
R4227 VSS.n1084 VSS 0.522821
R4228 VSS.n1050 VSS 0.522821
R4229 VSS.n1006 VSS 0.522821
R4230 VSS.n972 VSS 0.522821
R4231 VSS.n928 VSS 0.522821
R4232 VSS.n894 VSS 0.522821
R4233 VSS VSS.n1181 0.522821
R4234 VSS.n845 VSS.n844 0.517167
R4235 VSS.n1086 VSS.n853 0.517167
R4236 VSS.n1079 VSS.n1078 0.517167
R4237 VSS.n1045 VSS.n1044 0.517167
R4238 VSS.n1001 VSS.n1000 0.517167
R4239 VSS.n967 VSS.n966 0.517167
R4240 VSS.n923 VSS.n922 0.517167
R4241 VSS.n1180 VSS.n1179 0.517167
R4242 VSS.n847 VSS 0.455857
R4243 VSS VSS.n1083 0.455857
R4244 VSS VSS.n1049 0.455857
R4245 VSS VSS.n1005 0.455857
R4246 VSS VSS.n971 0.455857
R4247 VSS VSS.n927 0.455857
R4248 VSS VSS.n893 0.455857
R4249 VSS VSS.n571 0.426281
R4250 VSS.n808 VSS.n785 0.376971
R4251 VSS.n1099 VSS.n1098 0.376971
R4252 VSS.n1110 VSS.n1109 0.376971
R4253 VSS.n1121 VSS.n1120 0.376971
R4254 VSS.n1132 VSS.n1131 0.376971
R4255 VSS.n1143 VSS.n1142 0.376971
R4256 VSS.n1154 VSS.n1153 0.376971
R4257 VSS.n1165 VSS.n1164 0.376971
R4258 VSS.n811 VSS.n810 0.324029
R4259 VSS.n789 VSS.n788 0.324029
R4260 VSS.n792 VSS.n791 0.324029
R4261 VSS.n722 VSS.n721 0.324029
R4262 VSS.n715 VSS.n714 0.324029
R4263 VSS.n707 VSS.n706 0.324029
R4264 VSS.n700 VSS.n699 0.324029
R4265 VSS.n692 VSS.n691 0.324029
R4266 VSS.n685 VSS.n684 0.324029
R4267 VSS.n677 VSS.n676 0.324029
R4268 VSS.n670 VSS.n669 0.324029
R4269 VSS.n662 VSS.n661 0.324029
R4270 VSS.n655 VSS.n654 0.324029
R4271 VSS.n647 VSS.n646 0.324029
R4272 VSS.n640 VSS.n639 0.324029
R4273 VSS.n99 VSS.n98 0.324029
R4274 VSS.n120 VSS.n119 0.247896
R4275 VSS.n124 VSS.n120 0.247896
R4276 VSS.n126 VSS.n125 0.247896
R4277 VSS.n134 VSS.n129 0.247896
R4278 VSS.n614 VSS.n135 0.247896
R4279 VSS.n614 VSS.n613 0.247896
R4280 VSS.n612 VSS.n611 0.247896
R4281 VSS.n610 VSS.n609 0.247896
R4282 VSS.n608 VSS.n607 0.247896
R4283 VSS.n607 VSS.n142 0.247896
R4284 VSS.n146 VSS.n145 0.247896
R4285 VSS.n160 VSS.n155 0.247896
R4286 VSS.n598 VSS.n161 0.247896
R4287 VSS.n598 VSS.n597 0.247896
R4288 VSS.n596 VSS.n595 0.247896
R4289 VSS.n594 VSS.n593 0.247896
R4290 VSS.n592 VSS.n591 0.247896
R4291 VSS.n591 VSS.n168 0.247896
R4292 VSS.n172 VSS.n171 0.247896
R4293 VSS.n186 VSS.n181 0.247896
R4294 VSS.n582 VSS.n187 0.247896
R4295 VSS.n582 VSS.n581 0.247896
R4296 VSS.n580 VSS.n579 0.247896
R4297 VSS.n578 VSS.n577 0.247896
R4298 VSS.n576 VSS.n575 0.247896
R4299 VSS.n575 VSS.n194 0.247896
R4300 VSS.n572 VSS.n198 0.247896
R4301 VSS.n816 VSS.n815 0.247896
R4302 VSS.n822 VSS.n817 0.247896
R4303 VSS.n822 VSS.n821 0.247896
R4304 VSS.n820 VSS.n773 0.247896
R4305 VSS.n772 VSS.n771 0.247896
R4306 VSS.n770 VSS.n769 0.247896
R4307 VSS.n769 VSS.n760 0.247896
R4308 VSS.n759 VSS.n0 0.247896
R4309 VSS.n1243 VSS.n1242 0.247896
R4310 VSS.n1241 VSS.n1240 0.247896
R4311 VSS.n1240 VSS.n5 0.247896
R4312 VSS.n9 VSS.n8 0.247896
R4313 VSS.n19 VSS.n14 0.247896
R4314 VSS.n1229 VSS.n20 0.247896
R4315 VSS.n1229 VSS.n1228 0.247896
R4316 VSS.n1227 VSS.n1226 0.247896
R4317 VSS.n1225 VSS.n1224 0.247896
R4318 VSS.n1223 VSS.n1222 0.247896
R4319 VSS.n1222 VSS.n27 0.247896
R4320 VSS.n31 VSS.n30 0.247896
R4321 VSS.n41 VSS.n36 0.247896
R4322 VSS.n1211 VSS.n42 0.247896
R4323 VSS.n1211 VSS.n1210 0.247896
R4324 VSS.n1209 VSS.n1208 0.247896
R4325 VSS.n1207 VSS.n1206 0.247896
R4326 VSS.n1205 VSS.n1204 0.247896
R4327 VSS.n1204 VSS.n49 0.247896
R4328 VSS.n53 VSS.n52 0.247896
R4329 VSS.n63 VSS.n58 0.247896
R4330 VSS.n1193 VSS.n64 0.247896
R4331 VSS.n1193 VSS.n1192 0.247896
R4332 VSS.n1191 VSS.n1190 0.247896
R4333 VSS.n1189 VSS.n1188 0.247896
R4334 VSS.n1187 VSS.n1186 0.247896
R4335 VSS.n1186 VSS.n71 0.247896
R4336 VSS.n1183 VSS.n75 0.247896
R4337 VSS.n845 VSS.n734 0.246036
R4338 VSS.n853 VSS.n852 0.246036
R4339 VSS.n1080 VSS.n1079 0.246036
R4340 VSS.n1046 VSS.n1045 0.246036
R4341 VSS.n1002 VSS.n1001 0.246036
R4342 VSS.n968 VSS.n967 0.246036
R4343 VSS.n924 VSS.n923 0.246036
R4344 VSS.n1180 VSS.n79 0.246036
R4345 VSS.n812 VSS.n811 0.239471
R4346 VSS.n793 VSS.n792 0.239471
R4347 VSS.n716 VSS.n715 0.239471
R4348 VSS.n701 VSS.n700 0.239471
R4349 VSS.n686 VSS.n685 0.239471
R4350 VSS.n671 VSS.n670 0.239471
R4351 VSS.n656 VSS.n655 0.239471
R4352 VSS.n641 VSS.n640 0.239471
R4353 VSS.n794 VSS.n789 0.232118
R4354 VSS.n721 VSS.n717 0.232118
R4355 VSS.n706 VSS.n702 0.232118
R4356 VSS.n691 VSS.n687 0.232118
R4357 VSS.n676 VSS.n672 0.232118
R4358 VSS.n661 VSS.n657 0.232118
R4359 VSS.n646 VSS.n642 0.232118
R4360 VSS.n98 VSS.n94 0.232118
R4361 VSS.n119 VSS.n117 0.229667
R4362 VSS.n125 VSS.n124 0.229667
R4363 VSS.n135 VSS.n134 0.229667
R4364 VSS.n613 VSS.n612 0.229667
R4365 VSS.n609 VSS.n608 0.229667
R4366 VSS.n145 VSS.n142 0.229667
R4367 VSS.n161 VSS.n160 0.229667
R4368 VSS.n597 VSS.n596 0.229667
R4369 VSS.n593 VSS.n592 0.229667
R4370 VSS.n171 VSS.n168 0.229667
R4371 VSS.n187 VSS.n186 0.229667
R4372 VSS.n581 VSS.n580 0.229667
R4373 VSS.n577 VSS.n576 0.229667
R4374 VSS.n198 VSS.n194 0.229667
R4375 VSS.n817 VSS.n816 0.229667
R4376 VSS.n821 VSS.n820 0.229667
R4377 VSS.n771 VSS.n770 0.229667
R4378 VSS.n760 VSS.n759 0.229667
R4379 VSS.n1242 VSS.n1241 0.229667
R4380 VSS.n8 VSS.n5 0.229667
R4381 VSS.n20 VSS.n19 0.229667
R4382 VSS.n1228 VSS.n1227 0.229667
R4383 VSS.n1224 VSS.n1223 0.229667
R4384 VSS.n30 VSS.n27 0.229667
R4385 VSS.n42 VSS.n41 0.229667
R4386 VSS.n1210 VSS.n1209 0.229667
R4387 VSS.n1206 VSS.n1205 0.229667
R4388 VSS.n52 VSS.n49 0.229667
R4389 VSS.n64 VSS.n63 0.229667
R4390 VSS.n1192 VSS.n1191 0.229667
R4391 VSS.n1188 VSS.n1187 0.229667
R4392 VSS.n75 VSS.n71 0.229667
R4393 VSS.n571 VSS.n199 0.212219
R4394 VSS.n780 VSS.n779 0.196929
R4395 VSS.n779 VSS.n734 0.196929
R4396 VSS.n851 VSS.n850 0.196929
R4397 VSS.n852 VSS.n851 0.196929
R4398 VSS.n1082 VSS.n1081 0.196929
R4399 VSS.n1081 VSS.n1080 0.196929
R4400 VSS.n1048 VSS.n1047 0.196929
R4401 VSS.n1047 VSS.n1046 0.196929
R4402 VSS.n1004 VSS.n1003 0.196929
R4403 VSS.n1003 VSS.n1002 0.196929
R4404 VSS.n970 VSS.n969 0.196929
R4405 VSS.n969 VSS.n968 0.196929
R4406 VSS.n926 VSS.n925 0.196929
R4407 VSS.n925 VSS.n924 0.196929
R4408 VSS.n892 VSS.n891 0.196929
R4409 VSS.n891 VSS.n79 0.196929
R4410 VSS.n538 VSS.n199 0.189302
R4411 VSS.n542 VSS.n533 0.189302
R4412 VSS.n546 VSS.n544 0.189302
R4413 VSS.n530 VSS.n529 0.189302
R4414 VSS.n480 VSS.n478 0.189302
R4415 VSS.n495 VSS.n494 0.189302
R4416 VSS.n502 VSS.n497 0.189302
R4417 VSS.n505 VSS.n504 0.189302
R4418 VSS.n302 VSS.n297 0.189302
R4419 VSS.n306 VSS.n305 0.189302
R4420 VSS.n315 VSS.n290 0.189302
R4421 VSS.n319 VSS.n318 0.189302
R4422 VSS.n328 VSS.n283 0.189302
R4423 VSS.n332 VSS.n331 0.189302
R4424 VSS.n341 VSS.n276 0.189302
R4425 VSS.n345 VSS.n344 0.189302
R4426 VSS.n354 VSS.n269 0.189302
R4427 VSS.n358 VSS.n357 0.189302
R4428 VSS.n367 VSS.n262 0.189302
R4429 VSS.n371 VSS.n370 0.189302
R4430 VSS.n380 VSS.n255 0.189302
R4431 VSS.n384 VSS.n383 0.189302
R4432 VSS.n393 VSS.n248 0.189302
R4433 VSS.n397 VSS.n396 0.189302
R4434 VSS.n406 VSS.n241 0.189302
R4435 VSS.n410 VSS.n409 0.189302
R4436 VSS.n419 VSS.n234 0.189302
R4437 VSS.n423 VSS.n422 0.189302
R4438 VSS.n432 VSS.n227 0.189302
R4439 VSS.n436 VSS.n435 0.189302
R4440 VSS.n445 VSS.n220 0.189302
R4441 VSS.n449 VSS.n448 0.189302
R4442 VSS.n458 VSS.n213 0.189302
R4443 VSS.n464 VSS.n463 0.189302
R4444 VSS.n461 VSS.n208 0.189302
R4445 VSS.n205 VSS.n204 0.189302
R4446 VSS VSS.n76 0.172069
R4447 VSS VSS.n126 0.147635
R4448 VSS.n611 VSS 0.147635
R4449 VSS VSS.n146 0.147635
R4450 VSS.n595 VSS 0.147635
R4451 VSS VSS.n172 0.147635
R4452 VSS.n579 VSS 0.147635
R4453 VSS.n572 VSS 0.147635
R4454 VSS.n773 VSS 0.147635
R4455 VSS VSS.n0 0.147635
R4456 VSS VSS.n9 0.147635
R4457 VSS.n1226 VSS 0.147635
R4458 VSS VSS.n31 0.147635
R4459 VSS.n1208 VSS 0.147635
R4460 VSS VSS.n53 0.147635
R4461 VSS.n1190 VSS 0.147635
R4462 VSS.n1183 VSS 0.147635
R4463 VSS.n781 VSS.n780 0.146705
R4464 VSS.n850 VSS.n847 0.146705
R4465 VSS.n1083 VSS.n1082 0.146705
R4466 VSS.n1049 VSS.n1048 0.146705
R4467 VSS.n1005 VSS.n1004 0.146705
R4468 VSS.n971 VSS.n970 0.146705
R4469 VSS.n927 VSS.n926 0.146705
R4470 VSS.n893 VSS.n892 0.146705
R4471 VSS.n537 VSS.n533 0.13201
R4472 VSS.n544 VSS.n543 0.13201
R4473 VSS.n545 VSS.n530 0.13201
R4474 VSS.n528 VSS.n478 0.13201
R4475 VSS.n494 VSS.n493 0.13201
R4476 VSS.n497 VSS.n496 0.13201
R4477 VSS.n504 VSS.n503 0.13201
R4478 VSS.n507 VSS.n506 0.13201
R4479 VSS.n306 VSS.n303 0.13201
R4480 VSS.n304 VSS.n290 0.13201
R4481 VSS.n319 VSS.n316 0.13201
R4482 VSS.n317 VSS.n283 0.13201
R4483 VSS.n332 VSS.n329 0.13201
R4484 VSS.n330 VSS.n276 0.13201
R4485 VSS.n345 VSS.n342 0.13201
R4486 VSS.n343 VSS.n269 0.13201
R4487 VSS.n358 VSS.n355 0.13201
R4488 VSS.n356 VSS.n262 0.13201
R4489 VSS.n371 VSS.n368 0.13201
R4490 VSS.n369 VSS.n255 0.13201
R4491 VSS.n384 VSS.n381 0.13201
R4492 VSS.n382 VSS.n248 0.13201
R4493 VSS.n397 VSS.n394 0.13201
R4494 VSS.n395 VSS.n241 0.13201
R4495 VSS.n410 VSS.n407 0.13201
R4496 VSS.n408 VSS.n234 0.13201
R4497 VSS.n423 VSS.n420 0.13201
R4498 VSS.n421 VSS.n227 0.13201
R4499 VSS.n436 VSS.n433 0.13201
R4500 VSS.n434 VSS.n220 0.13201
R4501 VSS.n449 VSS.n446 0.13201
R4502 VSS.n447 VSS.n213 0.13201
R4503 VSS.n464 VSS.n459 0.13201
R4504 VSS.n462 VSS.n461 0.13201
R4505 VSS.n207 VSS.n205 0.13201
R4506 VSS.n570 VSS.n200 0.13201
R4507 VSS.n788 VSS.n784 0.124275
R4508 VSS.n723 VSS.n722 0.124275
R4509 VSS.n708 VSS.n707 0.124275
R4510 VSS.n693 VSS.n692 0.124275
R4511 VSS.n678 VSS.n677 0.124275
R4512 VSS.n663 VSS.n662 0.124275
R4513 VSS.n648 VSS.n647 0.124275
R4514 VSS.n100 VSS.n99 0.124275
R4515 VSS.n810 VSS.n809 0.120598
R4516 VSS.n791 VSS.n724 0.120598
R4517 VSS.n714 VSS.n709 0.120598
R4518 VSS.n699 VSS.n694 0.120598
R4519 VSS.n684 VSS.n679 0.120598
R4520 VSS.n669 VSS.n664 0.120598
R4521 VSS.n654 VSS.n649 0.120598
R4522 VSS.n639 VSS.n101 0.120598
R4523 VSS.n794 VSS 0.113245
R4524 VSS.n717 VSS 0.113245
R4525 VSS.n702 VSS 0.113245
R4526 VSS.n687 VSS 0.113245
R4527 VSS.n672 VSS 0.113245
R4528 VSS.n657 VSS 0.113245
R4529 VSS.n642 VSS 0.113245
R4530 VSS.n94 VSS 0.113245
R4531 VSS.n129 VSS 0.0721146
R4532 VSS VSS.n610 0.0721146
R4533 VSS.n155 VSS 0.0721146
R4534 VSS VSS.n594 0.0721146
R4535 VSS.n181 VSS 0.0721146
R4536 VSS VSS.n578 0.0721146
R4537 VSS.n507 VSS 0.0708125
R4538 VSS VSS.n570 0.0708125
R4539 VSS.n538 VSS.n537 0.0577917
R4540 VSS.n543 VSS.n542 0.0577917
R4541 VSS.n546 VSS.n545 0.0577917
R4542 VSS.n529 VSS.n528 0.0577917
R4543 VSS.n493 VSS.n480 0.0577917
R4544 VSS.n496 VSS.n495 0.0577917
R4545 VSS.n503 VSS.n502 0.0577917
R4546 VSS.n506 VSS.n505 0.0577917
R4547 VSS.n303 VSS.n302 0.0577917
R4548 VSS.n305 VSS.n304 0.0577917
R4549 VSS.n316 VSS.n315 0.0577917
R4550 VSS.n318 VSS.n317 0.0577917
R4551 VSS.n329 VSS.n328 0.0577917
R4552 VSS.n331 VSS.n330 0.0577917
R4553 VSS.n342 VSS.n341 0.0577917
R4554 VSS.n344 VSS.n343 0.0577917
R4555 VSS.n355 VSS.n354 0.0577917
R4556 VSS.n357 VSS.n356 0.0577917
R4557 VSS.n368 VSS.n367 0.0577917
R4558 VSS.n370 VSS.n369 0.0577917
R4559 VSS.n381 VSS.n380 0.0577917
R4560 VSS.n383 VSS.n382 0.0577917
R4561 VSS.n394 VSS.n393 0.0577917
R4562 VSS.n396 VSS.n395 0.0577917
R4563 VSS.n407 VSS.n406 0.0577917
R4564 VSS.n409 VSS.n408 0.0577917
R4565 VSS.n420 VSS.n419 0.0577917
R4566 VSS.n422 VSS.n421 0.0577917
R4567 VSS.n433 VSS.n432 0.0577917
R4568 VSS.n435 VSS.n434 0.0577917
R4569 VSS.n446 VSS.n445 0.0577917
R4570 VSS.n448 VSS.n447 0.0577917
R4571 VSS.n459 VSS.n458 0.0577917
R4572 VSS.n463 VSS.n462 0.0577917
R4573 VSS.n208 VSS.n207 0.0577917
R4574 VSS.n204 VSS.n200 0.0577917
R4575 VSS.n809 VSS.n784 0.00417647
R4576 VSS.n724 VSS.n723 0.00417647
R4577 VSS.n709 VSS.n708 0.00417647
R4578 VSS.n694 VSS.n693 0.00417647
R4579 VSS.n679 VSS.n678 0.00417647
R4580 VSS.n664 VSS.n663 0.00417647
R4581 VSS.n649 VSS.n648 0.00417647
R4582 VSS.n101 VSS.n100 0.00417647
R4583 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 572.12
R4584 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 572.12
R4585 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 572.12
R4586 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 572.12
R4587 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 539.841
R4588 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 539.841
R4589 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 539.841
R4590 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 539.841
R4591 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 215.293
R4592 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 215.293
R4593 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 215.293
R4594 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 215.293
R4595 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 166.468
R4596 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 166.149
R4597 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 165.8
R4598 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 165.8
R4599 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 85.1574
R4600 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 83.8097
R4601 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 83.8097
R4602 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 83.7172
R4603 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 74.288
R4604 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 67.7574
R4605 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 36.1505
R4606 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 36.1505
R4607 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 34.5438
R4608 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 34.5438
R4609 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 17.4005
R4610 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 17.4005
R4611 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 16.0275
R4612 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 11.8364
R4613 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 9.52217
R4614 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 9.52217
R4615 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 6.02878
R4616 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 5.83219
R4617 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 5.74235
R4618 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 5.49235
R4619 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 1.44072
R4620 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 1.32081
R4621 a_14774_2192.t10 a_14774_2192.n10 32.0282
R4622 a_14774_2192.n5 a_14774_2192.n4 25.7663
R4623 a_14774_2192.n8 a_14774_2192.n2 25.75
R4624 a_14774_2192.n9 a_14774_2192.n1 25.75
R4625 a_14774_2192.n10 a_14774_2192.n0 25.75
R4626 a_14774_2192.n5 a_14774_2192.n3 25.288
R4627 a_14774_2192.n7 a_14774_2192.n6 24.288
R4628 a_14774_2192.n6 a_14774_2192.t12 5.8005
R4629 a_14774_2192.n6 a_14774_2192.t11 5.8005
R4630 a_14774_2192.n3 a_14774_2192.t1 5.8005
R4631 a_14774_2192.n3 a_14774_2192.t0 5.8005
R4632 a_14774_2192.n4 a_14774_2192.t5 5.8005
R4633 a_14774_2192.n4 a_14774_2192.t2 5.8005
R4634 a_14774_2192.n2 a_14774_2192.t4 5.8005
R4635 a_14774_2192.n2 a_14774_2192.t9 5.8005
R4636 a_14774_2192.n1 a_14774_2192.t7 5.8005
R4637 a_14774_2192.n1 a_14774_2192.t6 5.8005
R4638 a_14774_2192.n0 a_14774_2192.t3 5.8005
R4639 a_14774_2192.n0 a_14774_2192.t8 5.8005
R4640 a_14774_2192.n8 a_14774_2192.n7 1.94072
R4641 a_14774_2192.n7 a_14774_2192.n5 1.47876
R4642 a_14774_2192.n9 a_14774_2192.n8 0.478761
R4643 a_14774_2192.n10 a_14774_2192.n9 0.478761
R4644 diff_gen_0.delay_unit_2_5.in_2.n4 diff_gen_0.delay_unit_2_5.in_2.t14 539.841
R4645 diff_gen_0.delay_unit_2_5.in_2.n5 diff_gen_0.delay_unit_2_5.in_2.t9 539.841
R4646 diff_gen_0.delay_unit_2_5.in_2.n1 diff_gen_0.delay_unit_2_5.in_2.t13 539.841
R4647 diff_gen_0.delay_unit_2_5.in_2.n2 diff_gen_0.delay_unit_2_5.in_2.t10 539.841
R4648 diff_gen_0.delay_unit_2_5.in_2.n4 diff_gen_0.delay_unit_2_5.in_2.t8 215.293
R4649 diff_gen_0.delay_unit_2_5.in_2.n5 diff_gen_0.delay_unit_2_5.in_2.t11 215.293
R4650 diff_gen_0.delay_unit_2_5.in_2.n1 diff_gen_0.delay_unit_2_5.in_2.t15 215.293
R4651 diff_gen_0.delay_unit_2_5.in_2.n2 diff_gen_0.delay_unit_2_5.in_2.t12 215.293
R4652 diff_gen_0.delay_unit_2_5.in_2.n7 diff_gen_0.delay_unit_2_5.in_2.n3 166.144
R4653 diff_gen_0.delay_unit_2_5.in_2.n7 diff_gen_0.delay_unit_2_5.in_2.n6 165.8
R4654 diff_gen_0.delay_unit_2_5.in_2.n12 diff_gen_0.delay_unit_2_5.in_2.t3 85.2499
R4655 diff_gen_0.delay_unit_2_5.in_2.n8 diff_gen_0.delay_unit_2_5.in_2.t4 85.2499
R4656 diff_gen_0.delay_unit_2_5.in_2.n12 diff_gen_0.delay_unit_2_5.in_2.t5 83.7172
R4657 diff_gen_0.delay_unit_2_5.in_2.n8 diff_gen_0.delay_unit_2_5.in_2.t2 83.7172
R4658 diff_gen_0.delay_unit_2_5.in_2.n11 diff_gen_0.delay_unit_2_5.in_2.n9 75.7282
R4659 diff_gen_0.delay_unit_2_5.in_2.n11 diff_gen_0.delay_unit_2_5.in_2.n10 66.3172
R4660 diff_gen_0.delay_unit_2_5.in_2.n6 diff_gen_0.delay_unit_2_5.in_2.n4 36.1505
R4661 diff_gen_0.delay_unit_2_5.in_2.n3 diff_gen_0.delay_unit_2_5.in_2.n1 36.1505
R4662 diff_gen_0.delay_unit_2_5.in_2.n6 diff_gen_0.delay_unit_2_5.in_2.n5 34.5438
R4663 diff_gen_0.delay_unit_2_5.in_2.n3 diff_gen_0.delay_unit_2_5.in_2.n2 34.5438
R4664 diff_gen_0.delay_unit_2_5.in_2.n10 diff_gen_0.delay_unit_2_5.in_2.t6 17.4005
R4665 diff_gen_0.delay_unit_2_5.in_2.n10 diff_gen_0.delay_unit_2_5.in_2.t7 17.4005
R4666 diff_gen_0.delay_unit_2_5.in_2.n9 diff_gen_0.delay_unit_2_5.in_2.t0 9.52217
R4667 diff_gen_0.delay_unit_2_5.in_2.n9 diff_gen_0.delay_unit_2_5.in_2.t1 9.52217
R4668 diff_gen_0.delay_unit_2_5.in_2.n0 diff_gen_0.delay_unit_2_5.in_2.n8 6.45821
R4669 diff_gen_0.delay_unit_2_5.in_2.n0 diff_gen_0.delay_unit_2_5.in_2.n11 5.30824
R4670 diff_gen_0.delay_unit_2_5.in_2.n0 diff_gen_0.delay_unit_2_5.in_2.n12 4.94887
R4671 diff_gen_0.delay_unit_2_5.in_2.n0 diff_gen_0.delay_unit_2_5.in_2.n7 1.41456
R4672 diff_gen_0.delay_unit_2_6.in_1.n3 diff_gen_0.delay_unit_2_6.in_1.t14 539.841
R4673 diff_gen_0.delay_unit_2_6.in_1.n4 diff_gen_0.delay_unit_2_6.in_1.t12 539.841
R4674 diff_gen_0.delay_unit_2_6.in_1.n0 diff_gen_0.delay_unit_2_6.in_1.t13 539.841
R4675 diff_gen_0.delay_unit_2_6.in_1.n1 diff_gen_0.delay_unit_2_6.in_1.t10 539.841
R4676 diff_gen_0.delay_unit_2_6.in_1.n3 diff_gen_0.delay_unit_2_6.in_1.t9 215.293
R4677 diff_gen_0.delay_unit_2_6.in_1.n4 diff_gen_0.delay_unit_2_6.in_1.t15 215.293
R4678 diff_gen_0.delay_unit_2_6.in_1.n0 diff_gen_0.delay_unit_2_6.in_1.t8 215.293
R4679 diff_gen_0.delay_unit_2_6.in_1.n1 diff_gen_0.delay_unit_2_6.in_1.t11 215.293
R4680 diff_gen_0.delay_unit_2_6.in_1.n6 diff_gen_0.delay_unit_2_6.in_1.n2 166.149
R4681 diff_gen_0.delay_unit_2_6.in_1.n6 diff_gen_0.delay_unit_2_6.in_1.n5 165.8
R4682 diff_gen_0.delay_unit_2_6.in_1.n12 diff_gen_0.delay_unit_2_6.in_1.t0 85.1574
R4683 diff_gen_0.delay_unit_2_6.in_1.n7 diff_gen_0.delay_unit_2_6.in_1.t7 85.1574
R4684 diff_gen_0.delay_unit_2_6.in_1.n12 diff_gen_0.delay_unit_2_6.in_1.t4 83.8097
R4685 diff_gen_0.delay_unit_2_6.in_1.n7 diff_gen_0.delay_unit_2_6.in_1.t6 83.8097
R4686 diff_gen_0.delay_unit_2_6.in_1.n11 diff_gen_0.delay_unit_2_6.in_1.n10 74.288
R4687 diff_gen_0.delay_unit_2_6.in_1.n11 diff_gen_0.delay_unit_2_6.in_1.n9 67.7574
R4688 diff_gen_0.delay_unit_2_6.in_1.n5 diff_gen_0.delay_unit_2_6.in_1.n3 36.1505
R4689 diff_gen_0.delay_unit_2_6.in_1.n2 diff_gen_0.delay_unit_2_6.in_1.n1 36.1505
R4690 diff_gen_0.delay_unit_2_6.in_1.n5 diff_gen_0.delay_unit_2_6.in_1.n4 34.5438
R4691 diff_gen_0.delay_unit_2_6.in_1.n2 diff_gen_0.delay_unit_2_6.in_1.n0 34.5438
R4692 diff_gen_0.delay_unit_2_6.in_1.n9 diff_gen_0.delay_unit_2_6.in_1.t1 17.4005
R4693 diff_gen_0.delay_unit_2_6.in_1.n9 diff_gen_0.delay_unit_2_6.in_1.t2 17.4005
R4694 diff_gen_0.delay_unit_2_6.in_1.n8 diff_gen_0.delay_unit_2_6.in_1.n6 11.8364
R4695 diff_gen_0.delay_unit_2_6.in_1.n10 diff_gen_0.delay_unit_2_6.in_1.t5 9.52217
R4696 diff_gen_0.delay_unit_2_6.in_1.n10 diff_gen_0.delay_unit_2_6.in_1.t3 9.52217
R4697 diff_gen_0.delay_unit_2_6.in_1.n13 diff_gen_0.delay_unit_2_6.in_1.n11 5.83219
R4698 diff_gen_0.delay_unit_2_6.in_1.n8 diff_gen_0.delay_unit_2_6.in_1.n7 5.74235
R4699 diff_gen_0.delay_unit_2_6.in_1.n13 diff_gen_0.delay_unit_2_6.in_1.n12 5.49235
R4700 diff_gen_0.delay_unit_2_6.in_1 diff_gen_0.delay_unit_2_6.in_1.n13 1.32081
R4701 diff_gen_0.delay_unit_2_6.in_1 diff_gen_0.delay_unit_2_6.in_1.n8 0.285656
R4702 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 879.481
R4703 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 742.783
R4704 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 665.16
R4705 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 623.388
R4706 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 523.774
R4707 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 431.807
R4708 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 427.875
R4709 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 357.26
R4710 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 208.537
R4711 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 168.077
R4712 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R4713 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R4714 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 31.2347
R4715 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 11.1806
R4716 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R4717 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R4718 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R4719 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R4720 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R4721 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 879.481
R4722 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 742.783
R4723 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 665.16
R4724 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 623.388
R4725 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 523.774
R4726 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 431.807
R4727 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 427.875
R4728 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 357.26
R4729 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 208.537
R4730 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 168.077
R4731 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R4732 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R4733 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 31.2347
R4734 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 11.1806
R4735 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R4736 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R4737 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R4738 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R4739 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R4740 vernier_delay_line_0.stop_strong.n0 vernier_delay_line_0.stop_strong.t79 851.506
R4741 vernier_delay_line_0.stop_strong.n78 vernier_delay_line_0.stop_strong.t51 851.506
R4742 vernier_delay_line_0.stop_strong.n71 vernier_delay_line_0.stop_strong.t37 851.506
R4743 vernier_delay_line_0.stop_strong.n64 vernier_delay_line_0.stop_strong.t71 851.506
R4744 vernier_delay_line_0.stop_strong.n57 vernier_delay_line_0.stop_strong.t56 851.506
R4745 vernier_delay_line_0.stop_strong.n50 vernier_delay_line_0.stop_strong.t85 851.506
R4746 vernier_delay_line_0.stop_strong.n43 vernier_delay_line_0.stop_strong.t74 851.506
R4747 vernier_delay_line_0.stop_strong.n36 vernier_delay_line_0.stop_strong.t64 851.506
R4748 vernier_delay_line_0.stop_strong.n0 vernier_delay_line_0.stop_strong.t75 850.414
R4749 vernier_delay_line_0.stop_strong.n78 vernier_delay_line_0.stop_strong.t54 850.414
R4750 vernier_delay_line_0.stop_strong.n71 vernier_delay_line_0.stop_strong.t40 850.414
R4751 vernier_delay_line_0.stop_strong.n64 vernier_delay_line_0.stop_strong.t68 850.414
R4752 vernier_delay_line_0.stop_strong.n57 vernier_delay_line_0.stop_strong.t60 850.414
R4753 vernier_delay_line_0.stop_strong.n50 vernier_delay_line_0.stop_strong.t45 850.414
R4754 vernier_delay_line_0.stop_strong.n43 vernier_delay_line_0.stop_strong.t77 850.414
R4755 vernier_delay_line_0.stop_strong.n36 vernier_delay_line_0.stop_strong.t50 850.414
R4756 vernier_delay_line_0.stop_strong.n1 vernier_delay_line_0.stop_strong.t80 665.16
R4757 vernier_delay_line_0.stop_strong.n79 vernier_delay_line_0.stop_strong.t67 665.16
R4758 vernier_delay_line_0.stop_strong.n72 vernier_delay_line_0.stop_strong.t62 665.16
R4759 vernier_delay_line_0.stop_strong.n65 vernier_delay_line_0.stop_strong.t86 665.16
R4760 vernier_delay_line_0.stop_strong.n58 vernier_delay_line_0.stop_strong.t87 665.16
R4761 vernier_delay_line_0.stop_strong.n51 vernier_delay_line_0.stop_strong.t49 665.16
R4762 vernier_delay_line_0.stop_strong.n44 vernier_delay_line_0.stop_strong.t36 665.16
R4763 vernier_delay_line_0.stop_strong.n37 vernier_delay_line_0.stop_strong.t65 665.16
R4764 vernier_delay_line_0.stop_strong.n1 vernier_delay_line_0.stop_strong.t59 523.774
R4765 vernier_delay_line_0.stop_strong.n2 vernier_delay_line_0.stop_strong.t43 523.774
R4766 vernier_delay_line_0.stop_strong.n3 vernier_delay_line_0.stop_strong.t38 523.774
R4767 vernier_delay_line_0.stop_strong.n4 vernier_delay_line_0.stop_strong.t72 523.774
R4768 vernier_delay_line_0.stop_strong.n79 vernier_delay_line_0.stop_strong.t44 523.774
R4769 vernier_delay_line_0.stop_strong.n80 vernier_delay_line_0.stop_strong.t76 523.774
R4770 vernier_delay_line_0.stop_strong.n81 vernier_delay_line_0.stop_strong.t55 523.774
R4771 vernier_delay_line_0.stop_strong.n82 vernier_delay_line_0.stop_strong.t83 523.774
R4772 vernier_delay_line_0.stop_strong.n72 vernier_delay_line_0.stop_strong.t32 523.774
R4773 vernier_delay_line_0.stop_strong.n73 vernier_delay_line_0.stop_strong.t66 523.774
R4774 vernier_delay_line_0.stop_strong.n74 vernier_delay_line_0.stop_strong.t84 523.774
R4775 vernier_delay_line_0.stop_strong.n75 vernier_delay_line_0.stop_strong.t63 523.774
R4776 vernier_delay_line_0.stop_strong.n65 vernier_delay_line_0.stop_strong.t82 523.774
R4777 vernier_delay_line_0.stop_strong.n66 vernier_delay_line_0.stop_strong.t41 523.774
R4778 vernier_delay_line_0.stop_strong.n67 vernier_delay_line_0.stop_strong.t73 523.774
R4779 vernier_delay_line_0.stop_strong.n68 vernier_delay_line_0.stop_strong.t52 523.774
R4780 vernier_delay_line_0.stop_strong.n58 vernier_delay_line_0.stop_strong.t48 523.774
R4781 vernier_delay_line_0.stop_strong.n59 vernier_delay_line_0.stop_strong.t81 523.774
R4782 vernier_delay_line_0.stop_strong.n60 vernier_delay_line_0.stop_strong.t61 523.774
R4783 vernier_delay_line_0.stop_strong.n61 vernier_delay_line_0.stop_strong.t53 523.774
R4784 vernier_delay_line_0.stop_strong.n51 vernier_delay_line_0.stop_strong.t35 523.774
R4785 vernier_delay_line_0.stop_strong.n52 vernier_delay_line_0.stop_strong.t69 523.774
R4786 vernier_delay_line_0.stop_strong.n53 vernier_delay_line_0.stop_strong.t46 523.774
R4787 vernier_delay_line_0.stop_strong.n54 vernier_delay_line_0.stop_strong.t78 523.774
R4788 vernier_delay_line_0.stop_strong.n44 vernier_delay_line_0.stop_strong.t70 523.774
R4789 vernier_delay_line_0.stop_strong.n45 vernier_delay_line_0.stop_strong.t47 523.774
R4790 vernier_delay_line_0.stop_strong.n46 vernier_delay_line_0.stop_strong.t33 523.774
R4791 vernier_delay_line_0.stop_strong.n47 vernier_delay_line_0.stop_strong.t57 523.774
R4792 vernier_delay_line_0.stop_strong.n37 vernier_delay_line_0.stop_strong.t39 523.774
R4793 vernier_delay_line_0.stop_strong.n38 vernier_delay_line_0.stop_strong.t34 523.774
R4794 vernier_delay_line_0.stop_strong.n39 vernier_delay_line_0.stop_strong.t58 523.774
R4795 vernier_delay_line_0.stop_strong.n40 vernier_delay_line_0.stop_strong.t42 523.774
R4796 vernier_delay_line_0.stop_strong.n5 vernier_delay_line_0.stop_strong.n4 213.51
R4797 vernier_delay_line_0.stop_strong.n83 vernier_delay_line_0.stop_strong.n82 213.51
R4798 vernier_delay_line_0.stop_strong.n76 vernier_delay_line_0.stop_strong.n75 213.51
R4799 vernier_delay_line_0.stop_strong.n69 vernier_delay_line_0.stop_strong.n68 213.51
R4800 vernier_delay_line_0.stop_strong.n62 vernier_delay_line_0.stop_strong.n61 213.51
R4801 vernier_delay_line_0.stop_strong.n55 vernier_delay_line_0.stop_strong.n54 213.51
R4802 vernier_delay_line_0.stop_strong.n48 vernier_delay_line_0.stop_strong.n47 213.51
R4803 vernier_delay_line_0.stop_strong.n41 vernier_delay_line_0.stop_strong.n40 213.51
R4804 vernier_delay_line_0.stop_strong.n4 vernier_delay_line_0.stop_strong.n3 141.387
R4805 vernier_delay_line_0.stop_strong.n3 vernier_delay_line_0.stop_strong.n2 141.387
R4806 vernier_delay_line_0.stop_strong.n2 vernier_delay_line_0.stop_strong.n1 141.387
R4807 vernier_delay_line_0.stop_strong.n82 vernier_delay_line_0.stop_strong.n81 141.387
R4808 vernier_delay_line_0.stop_strong.n81 vernier_delay_line_0.stop_strong.n80 141.387
R4809 vernier_delay_line_0.stop_strong.n80 vernier_delay_line_0.stop_strong.n79 141.387
R4810 vernier_delay_line_0.stop_strong.n75 vernier_delay_line_0.stop_strong.n74 141.387
R4811 vernier_delay_line_0.stop_strong.n74 vernier_delay_line_0.stop_strong.n73 141.387
R4812 vernier_delay_line_0.stop_strong.n73 vernier_delay_line_0.stop_strong.n72 141.387
R4813 vernier_delay_line_0.stop_strong.n68 vernier_delay_line_0.stop_strong.n67 141.387
R4814 vernier_delay_line_0.stop_strong.n67 vernier_delay_line_0.stop_strong.n66 141.387
R4815 vernier_delay_line_0.stop_strong.n66 vernier_delay_line_0.stop_strong.n65 141.387
R4816 vernier_delay_line_0.stop_strong.n61 vernier_delay_line_0.stop_strong.n60 141.387
R4817 vernier_delay_line_0.stop_strong.n60 vernier_delay_line_0.stop_strong.n59 141.387
R4818 vernier_delay_line_0.stop_strong.n59 vernier_delay_line_0.stop_strong.n58 141.387
R4819 vernier_delay_line_0.stop_strong.n54 vernier_delay_line_0.stop_strong.n53 141.387
R4820 vernier_delay_line_0.stop_strong.n53 vernier_delay_line_0.stop_strong.n52 141.387
R4821 vernier_delay_line_0.stop_strong.n52 vernier_delay_line_0.stop_strong.n51 141.387
R4822 vernier_delay_line_0.stop_strong.n47 vernier_delay_line_0.stop_strong.n46 141.387
R4823 vernier_delay_line_0.stop_strong.n46 vernier_delay_line_0.stop_strong.n45 141.387
R4824 vernier_delay_line_0.stop_strong.n45 vernier_delay_line_0.stop_strong.n44 141.387
R4825 vernier_delay_line_0.stop_strong.n40 vernier_delay_line_0.stop_strong.n39 141.387
R4826 vernier_delay_line_0.stop_strong.n39 vernier_delay_line_0.stop_strong.n38 141.387
R4827 vernier_delay_line_0.stop_strong.n38 vernier_delay_line_0.stop_strong.n37 141.387
R4828 vernier_delay_line_0.stop_strong.n6 vernier_delay_line_0.stop_strong.t21 85.2499
R4829 vernier_delay_line_0.stop_strong.n7 vernier_delay_line_0.stop_strong.t9 85.2499
R4830 vernier_delay_line_0.stop_strong.n9 vernier_delay_line_0.stop_strong.t3 85.2499
R4831 vernier_delay_line_0.stop_strong.n11 vernier_delay_line_0.stop_strong.t18 85.2499
R4832 vernier_delay_line_0.stop_strong.n13 vernier_delay_line_0.stop_strong.t6 85.2499
R4833 vernier_delay_line_0.stop_strong.n15 vernier_delay_line_0.stop_strong.t15 85.2499
R4834 vernier_delay_line_0.stop_strong.n19 vernier_delay_line_0.stop_strong.t10 85.2499
R4835 vernier_delay_line_0.stop_strong.n21 vernier_delay_line_0.stop_strong.t31 85.2499
R4836 vernier_delay_line_0.stop_strong.n23 vernier_delay_line_0.stop_strong.t24 85.2499
R4837 vernier_delay_line_0.stop_strong.n25 vernier_delay_line_0.stop_strong.t13 85.2499
R4838 vernier_delay_line_0.stop_strong.n27 vernier_delay_line_0.stop_strong.t5 85.2499
R4839 vernier_delay_line_0.stop_strong.n29 vernier_delay_line_0.stop_strong.t23 85.2499
R4840 vernier_delay_line_0.stop_strong.n31 vernier_delay_line_0.stop_strong.t19 85.2499
R4841 vernier_delay_line_0.stop_strong.n33 vernier_delay_line_0.stop_strong.t7 85.2499
R4842 vernier_delay_line_0.stop_strong.n17 vernier_delay_line_0.stop_strong.t0 85.2499
R4843 stop_buffer_0.stop_strong vernier_delay_line_0.stop_strong.t26 84.7281
R4844 vernier_delay_line_0.stop_strong.n17 vernier_delay_line_0.stop_strong.t1 83.7172
R4845 vernier_delay_line_0.stop_strong.n6 vernier_delay_line_0.stop_strong.t16 83.7172
R4846 vernier_delay_line_0.stop_strong.n7 vernier_delay_line_0.stop_strong.t14 83.7172
R4847 vernier_delay_line_0.stop_strong.n9 vernier_delay_line_0.stop_strong.t28 83.7172
R4848 vernier_delay_line_0.stop_strong.n11 vernier_delay_line_0.stop_strong.t20 83.7172
R4849 vernier_delay_line_0.stop_strong.n13 vernier_delay_line_0.stop_strong.t8 83.7172
R4850 vernier_delay_line_0.stop_strong.n15 vernier_delay_line_0.stop_strong.t2 83.7172
R4851 vernier_delay_line_0.stop_strong.n19 vernier_delay_line_0.stop_strong.t11 83.7172
R4852 vernier_delay_line_0.stop_strong.n21 vernier_delay_line_0.stop_strong.t22 83.7172
R4853 vernier_delay_line_0.stop_strong.n23 vernier_delay_line_0.stop_strong.t25 83.7172
R4854 vernier_delay_line_0.stop_strong.n25 vernier_delay_line_0.stop_strong.t17 83.7172
R4855 vernier_delay_line_0.stop_strong.n27 vernier_delay_line_0.stop_strong.t30 83.7172
R4856 vernier_delay_line_0.stop_strong.n29 vernier_delay_line_0.stop_strong.t29 83.7172
R4857 vernier_delay_line_0.stop_strong.n31 vernier_delay_line_0.stop_strong.t12 83.7172
R4858 vernier_delay_line_0.stop_strong.n33 vernier_delay_line_0.stop_strong.t4 83.7172
R4859 stop_buffer_0.stop_strong vernier_delay_line_0.stop_strong.t27 83.7172
R4860 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n5 11.8482
R4861 vernier_delay_line_0.stop_strong.n84 vernier_delay_line_0.stop_strong.n83 9.66066
R4862 vernier_delay_line_0.stop_strong.n77 vernier_delay_line_0.stop_strong.n76 9.66066
R4863 vernier_delay_line_0.stop_strong.n70 vernier_delay_line_0.stop_strong.n69 9.66066
R4864 vernier_delay_line_0.stop_strong.n63 vernier_delay_line_0.stop_strong.n62 9.66066
R4865 vernier_delay_line_0.stop_strong.n56 vernier_delay_line_0.stop_strong.n55 9.66066
R4866 vernier_delay_line_0.stop_strong.n49 vernier_delay_line_0.stop_strong.n48 9.66066
R4867 vernier_delay_line_0.stop_strong.n42 vernier_delay_line_0.stop_strong.n41 9.66066
R4868 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n35 8.04701
R4869 vernier_delay_line_0.stop_strong.n8 vernier_delay_line_0.stop_strong.n6 5.16238
R4870 vernier_delay_line_0.stop_strong.n35 stop_buffer_0.stop_strong 5.01952
R4871 vernier_delay_line_0.stop_strong.n8 vernier_delay_line_0.stop_strong.n7 4.64452
R4872 vernier_delay_line_0.stop_strong.n10 vernier_delay_line_0.stop_strong.n9 4.64452
R4873 vernier_delay_line_0.stop_strong.n12 vernier_delay_line_0.stop_strong.n11 4.64452
R4874 vernier_delay_line_0.stop_strong.n14 vernier_delay_line_0.stop_strong.n13 4.64452
R4875 vernier_delay_line_0.stop_strong.n16 vernier_delay_line_0.stop_strong.n15 4.64452
R4876 vernier_delay_line_0.stop_strong.n20 vernier_delay_line_0.stop_strong.n19 4.64452
R4877 vernier_delay_line_0.stop_strong.n22 vernier_delay_line_0.stop_strong.n21 4.64452
R4878 vernier_delay_line_0.stop_strong.n24 vernier_delay_line_0.stop_strong.n23 4.64452
R4879 vernier_delay_line_0.stop_strong.n26 vernier_delay_line_0.stop_strong.n25 4.64452
R4880 vernier_delay_line_0.stop_strong.n28 vernier_delay_line_0.stop_strong.n27 4.64452
R4881 vernier_delay_line_0.stop_strong.n30 vernier_delay_line_0.stop_strong.n29 4.64452
R4882 vernier_delay_line_0.stop_strong.n32 vernier_delay_line_0.stop_strong.n31 4.64452
R4883 vernier_delay_line_0.stop_strong.n34 vernier_delay_line_0.stop_strong.n33 4.64452
R4884 vernier_delay_line_0.stop_strong.n18 vernier_delay_line_0.stop_strong.n17 4.64452
R4885 vernier_delay_line_0.stop_strong.n84 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk 2.188
R4886 vernier_delay_line_0.stop_strong.n77 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk 2.188
R4887 vernier_delay_line_0.stop_strong.n70 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk 2.188
R4888 vernier_delay_line_0.stop_strong.n63 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk 2.188
R4889 vernier_delay_line_0.stop_strong.n56 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk 2.188
R4890 vernier_delay_line_0.stop_strong.n49 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk 2.188
R4891 vernier_delay_line_0.stop_strong.n42 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk 2.188
R4892 vernier_delay_line_0.stop_strong.n5 vernier_delay_line_0.stop_strong.n0 1.05649
R4893 vernier_delay_line_0.stop_strong.n83 vernier_delay_line_0.stop_strong.n78 1.05649
R4894 vernier_delay_line_0.stop_strong.n76 vernier_delay_line_0.stop_strong.n71 1.05649
R4895 vernier_delay_line_0.stop_strong.n69 vernier_delay_line_0.stop_strong.n64 1.05649
R4896 vernier_delay_line_0.stop_strong.n62 vernier_delay_line_0.stop_strong.n57 1.05649
R4897 vernier_delay_line_0.stop_strong.n55 vernier_delay_line_0.stop_strong.n50 1.05649
R4898 vernier_delay_line_0.stop_strong.n48 vernier_delay_line_0.stop_strong.n43 1.05649
R4899 vernier_delay_line_0.stop_strong.n41 vernier_delay_line_0.stop_strong.n36 1.05649
R4900 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n84 0.6655
R4901 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n77 0.6655
R4902 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n70 0.6655
R4903 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n63 0.6655
R4904 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n56 0.6655
R4905 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n49 0.6655
R4906 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk vernier_delay_line_0.stop_strong.n42 0.6655
R4907 vernier_delay_line_0.stop_strong.n34 vernier_delay_line_0.stop_strong.n32 0.518357
R4908 vernier_delay_line_0.stop_strong.n32 vernier_delay_line_0.stop_strong.n30 0.518357
R4909 vernier_delay_line_0.stop_strong.n30 vernier_delay_line_0.stop_strong.n28 0.518357
R4910 vernier_delay_line_0.stop_strong.n28 vernier_delay_line_0.stop_strong.n26 0.518357
R4911 vernier_delay_line_0.stop_strong.n26 vernier_delay_line_0.stop_strong.n24 0.518357
R4912 vernier_delay_line_0.stop_strong.n24 vernier_delay_line_0.stop_strong.n22 0.518357
R4913 vernier_delay_line_0.stop_strong.n22 vernier_delay_line_0.stop_strong.n20 0.518357
R4914 vernier_delay_line_0.stop_strong.n20 vernier_delay_line_0.stop_strong.n18 0.518357
R4915 vernier_delay_line_0.stop_strong.n18 vernier_delay_line_0.stop_strong.n16 0.518357
R4916 vernier_delay_line_0.stop_strong.n16 vernier_delay_line_0.stop_strong.n14 0.518357
R4917 vernier_delay_line_0.stop_strong.n14 vernier_delay_line_0.stop_strong.n12 0.518357
R4918 vernier_delay_line_0.stop_strong.n12 vernier_delay_line_0.stop_strong.n10 0.518357
R4919 vernier_delay_line_0.stop_strong.n10 vernier_delay_line_0.stop_strong.n8 0.518357
R4920 vernier_delay_line_0.stop_strong.n35 vernier_delay_line_0.stop_strong.n34 0.497131
R4921 a_12492_2192.n4 a_12492_2192.t10 32.0282
R4922 a_12492_2192.n9 a_12492_2192.n0 25.7663
R4923 a_12492_2192.n6 a_12492_2192.n1 25.75
R4924 a_12492_2192.n5 a_12492_2192.n2 25.75
R4925 a_12492_2192.n4 a_12492_2192.n3 25.75
R4926 a_12492_2192.n10 a_12492_2192.n9 25.288
R4927 a_12492_2192.n8 a_12492_2192.n7 24.288
R4928 a_12492_2192.n7 a_12492_2192.t8 5.8005
R4929 a_12492_2192.n7 a_12492_2192.t11 5.8005
R4930 a_12492_2192.n1 a_12492_2192.t12 5.8005
R4931 a_12492_2192.n1 a_12492_2192.t3 5.8005
R4932 a_12492_2192.n2 a_12492_2192.t2 5.8005
R4933 a_12492_2192.n2 a_12492_2192.t1 5.8005
R4934 a_12492_2192.n3 a_12492_2192.t4 5.8005
R4935 a_12492_2192.n3 a_12492_2192.t0 5.8005
R4936 a_12492_2192.n0 a_12492_2192.t7 5.8005
R4937 a_12492_2192.n0 a_12492_2192.t5 5.8005
R4938 a_12492_2192.n10 a_12492_2192.t6 5.8005
R4939 a_12492_2192.t9 a_12492_2192.n10 5.8005
R4940 a_12492_2192.n8 a_12492_2192.n6 1.94072
R4941 a_12492_2192.n9 a_12492_2192.n8 1.47876
R4942 a_12492_2192.n6 a_12492_2192.n5 0.478761
R4943 a_12492_2192.n5 a_12492_2192.n4 0.478761
R4944 diff_gen_0.delay_unit_2_2.in_1.n3 diff_gen_0.delay_unit_2_2.in_1.t11 539.841
R4945 diff_gen_0.delay_unit_2_2.in_1.n4 diff_gen_0.delay_unit_2_2.in_1.t10 539.841
R4946 diff_gen_0.delay_unit_2_2.in_1.n0 diff_gen_0.delay_unit_2_2.in_1.t9 539.841
R4947 diff_gen_0.delay_unit_2_2.in_1.n1 diff_gen_0.delay_unit_2_2.in_1.t15 539.841
R4948 diff_gen_0.delay_unit_2_2.in_1.n3 diff_gen_0.delay_unit_2_2.in_1.t14 215.293
R4949 diff_gen_0.delay_unit_2_2.in_1.n4 diff_gen_0.delay_unit_2_2.in_1.t13 215.293
R4950 diff_gen_0.delay_unit_2_2.in_1.n0 diff_gen_0.delay_unit_2_2.in_1.t12 215.293
R4951 diff_gen_0.delay_unit_2_2.in_1.n1 diff_gen_0.delay_unit_2_2.in_1.t8 215.293
R4952 diff_gen_0.delay_unit_2_2.in_1.n6 diff_gen_0.delay_unit_2_2.in_1.n2 166.149
R4953 diff_gen_0.delay_unit_2_2.in_1.n6 diff_gen_0.delay_unit_2_2.in_1.n5 165.8
R4954 diff_gen_0.delay_unit_2_2.in_1.n12 diff_gen_0.delay_unit_2_2.in_1.t7 85.1574
R4955 diff_gen_0.delay_unit_2_2.in_1.n7 diff_gen_0.delay_unit_2_2.in_1.t6 85.1574
R4956 diff_gen_0.delay_unit_2_2.in_1.n7 diff_gen_0.delay_unit_2_2.in_1.t4 83.8097
R4957 diff_gen_0.delay_unit_2_2.in_1.n12 diff_gen_0.delay_unit_2_2.in_1.t1 83.8097
R4958 diff_gen_0.delay_unit_2_2.in_1.n11 diff_gen_0.delay_unit_2_2.in_1.n10 74.288
R4959 diff_gen_0.delay_unit_2_2.in_1.n11 diff_gen_0.delay_unit_2_2.in_1.n9 67.7574
R4960 diff_gen_0.delay_unit_2_2.in_1.n5 diff_gen_0.delay_unit_2_2.in_1.n3 36.1505
R4961 diff_gen_0.delay_unit_2_2.in_1.n2 diff_gen_0.delay_unit_2_2.in_1.n1 36.1505
R4962 diff_gen_0.delay_unit_2_2.in_1.n5 diff_gen_0.delay_unit_2_2.in_1.n4 34.5438
R4963 diff_gen_0.delay_unit_2_2.in_1.n2 diff_gen_0.delay_unit_2_2.in_1.n0 34.5438
R4964 diff_gen_0.delay_unit_2_2.in_1.n9 diff_gen_0.delay_unit_2_2.in_1.t5 17.4005
R4965 diff_gen_0.delay_unit_2_2.in_1.n9 diff_gen_0.delay_unit_2_2.in_1.t0 17.4005
R4966 diff_gen_0.delay_unit_2_2.in_1.n8 diff_gen_0.delay_unit_2_2.in_1.n6 11.8364
R4967 diff_gen_0.delay_unit_2_2.in_1.n10 diff_gen_0.delay_unit_2_2.in_1.t3 9.52217
R4968 diff_gen_0.delay_unit_2_2.in_1.n10 diff_gen_0.delay_unit_2_2.in_1.t2 9.52217
R4969 diff_gen_0.delay_unit_2_2.in_1.n13 diff_gen_0.delay_unit_2_2.in_1.n11 5.83219
R4970 diff_gen_0.delay_unit_2_2.in_1.n8 diff_gen_0.delay_unit_2_2.in_1.n7 5.74235
R4971 diff_gen_0.delay_unit_2_2.in_1.n13 diff_gen_0.delay_unit_2_2.in_1.n12 5.49235
R4972 diff_gen_0.delay_unit_2_1.out_1 diff_gen_0.delay_unit_2_2.in_1.n13 1.32081
R4973 diff_gen_0.delay_unit_2_1.out_1 diff_gen_0.delay_unit_2_2.in_1.n8 0.53175
R4974 diff_gen_0.delay_unit_2_3.in_2.n3 diff_gen_0.delay_unit_2_3.in_2.t13 539.841
R4975 diff_gen_0.delay_unit_2_3.in_2.n4 diff_gen_0.delay_unit_2_3.in_2.t9 539.841
R4976 diff_gen_0.delay_unit_2_3.in_2.n0 diff_gen_0.delay_unit_2_3.in_2.t12 539.841
R4977 diff_gen_0.delay_unit_2_3.in_2.n1 diff_gen_0.delay_unit_2_3.in_2.t8 539.841
R4978 diff_gen_0.delay_unit_2_3.in_2.n3 diff_gen_0.delay_unit_2_3.in_2.t15 215.293
R4979 diff_gen_0.delay_unit_2_3.in_2.n4 diff_gen_0.delay_unit_2_3.in_2.t11 215.293
R4980 diff_gen_0.delay_unit_2_3.in_2.n0 diff_gen_0.delay_unit_2_3.in_2.t14 215.293
R4981 diff_gen_0.delay_unit_2_3.in_2.n1 diff_gen_0.delay_unit_2_3.in_2.t10 215.293
R4982 diff_gen_0.delay_unit_2_3.in_2.n6 diff_gen_0.delay_unit_2_3.in_2.n2 166.144
R4983 diff_gen_0.delay_unit_2_3.in_2.n6 diff_gen_0.delay_unit_2_3.in_2.n5 165.8
R4984 diff_gen_0.delay_unit_2_3.in_2.n7 diff_gen_0.delay_unit_2_3.in_2.t7 85.2499
R4985 diff_gen_0.delay_unit_2_3.in_2.n12 diff_gen_0.delay_unit_2_3.in_2.t5 85.2499
R4986 diff_gen_0.delay_unit_2_3.in_2.n12 diff_gen_0.delay_unit_2_3.in_2.t1 83.7172
R4987 diff_gen_0.delay_unit_2_3.in_2.n7 diff_gen_0.delay_unit_2_3.in_2.t6 83.7172
R4988 diff_gen_0.delay_unit_2_3.in_2.n11 diff_gen_0.delay_unit_2_3.in_2.n9 75.7282
R4989 diff_gen_0.delay_unit_2_3.in_2.n11 diff_gen_0.delay_unit_2_3.in_2.n10 66.3172
R4990 diff_gen_0.delay_unit_2_3.in_2.n5 diff_gen_0.delay_unit_2_3.in_2.n3 36.1505
R4991 diff_gen_0.delay_unit_2_3.in_2.n2 diff_gen_0.delay_unit_2_3.in_2.n0 36.1505
R4992 diff_gen_0.delay_unit_2_3.in_2.n5 diff_gen_0.delay_unit_2_3.in_2.n4 34.5438
R4993 diff_gen_0.delay_unit_2_3.in_2.n2 diff_gen_0.delay_unit_2_3.in_2.n1 34.5438
R4994 diff_gen_0.delay_unit_2_3.in_2.n10 diff_gen_0.delay_unit_2_3.in_2.t2 17.4005
R4995 diff_gen_0.delay_unit_2_3.in_2.n10 diff_gen_0.delay_unit_2_3.in_2.t0 17.4005
R4996 diff_gen_0.delay_unit_2_3.in_2.n9 diff_gen_0.delay_unit_2_3.in_2.t3 9.52217
R4997 diff_gen_0.delay_unit_2_3.in_2.n9 diff_gen_0.delay_unit_2_3.in_2.t4 9.52217
R4998 diff_gen_0.delay_unit_2_3.in_2.n8 diff_gen_0.delay_unit_2_3.in_2.n7 6.45821
R4999 diff_gen_0.delay_unit_2_3.in_2.n13 diff_gen_0.delay_unit_2_3.in_2.n11 5.30824
R5000 diff_gen_0.delay_unit_2_3.in_2.n13 diff_gen_0.delay_unit_2_3.in_2.n12 4.94887
R5001 diff_gen_0.delay_unit_2_3.in_2.n8 diff_gen_0.delay_unit_2_3.in_2.n6 1.06691
R5002 diff_gen_0.delay_unit_2_2.out_2 diff_gen_0.delay_unit_2_3.in_2.n8 0.188
R5003 diff_gen_0.delay_unit_2_2.out_2 diff_gen_0.delay_unit_2_3.in_2.n13 0.160656
R5004 start_buffer_0.start_buff.n12 start_buffer_0.start_buff.t19 543.053
R5005 start_buffer_0.start_buff.n11 start_buffer_0.start_buff.t22 543.053
R5006 start_buffer_0.start_buff.n10 start_buffer_0.start_buff.t15 543.053
R5007 start_buffer_0.start_buff.n3 start_buffer_0.start_buff.t17 539.841
R5008 start_buffer_0.start_buff.n4 start_buffer_0.start_buff.t10 539.841
R5009 start_buffer_0.start_buff.n0 start_buffer_0.start_buff.t11 539.841
R5010 start_buffer_0.start_buff.n1 start_buffer_0.start_buff.t21 539.841
R5011 start_buffer_0.start_buff.n12 start_buffer_0.start_buff.t20 221.72
R5012 start_buffer_0.start_buff.n11 start_buffer_0.start_buff.t23 221.72
R5013 start_buffer_0.start_buff.n10 start_buffer_0.start_buff.t16 221.72
R5014 start_buffer_0.start_buff.n13 start_buffer_0.start_buff.n11 218.32
R5015 start_buffer_0.start_buff.n13 start_buffer_0.start_buff.n12 217.734
R5016 start_buffer_0.start_buff.n3 start_buffer_0.start_buff.t18 215.293
R5017 start_buffer_0.start_buff.n4 start_buffer_0.start_buff.t13 215.293
R5018 start_buffer_0.start_buff.n0 start_buffer_0.start_buff.t14 215.293
R5019 start_buffer_0.start_buff.n1 start_buffer_0.start_buff.t12 215.293
R5020 start_buffer_0.start_buff.n14 start_buffer_0.start_buff.n10 213.234
R5021 start_buffer_0.start_buff.n6 start_buffer_0.start_buff.n2 166.149
R5022 start_buffer_0.start_buff.n6 start_buffer_0.start_buff.n5 165.8
R5023 start_buffer_0.start_buff.n17 start_buffer_0.start_buff.t4 85.2499
R5024 start_buffer_0.start_buff.n20 start_buffer_0.start_buff.t6 85.2499
R5025 start_buffer_0.start_buff.n18 start_buffer_0.start_buff.t7 85.2499
R5026 start_buffer_0.start_buff.n7 start_buffer_0.start_buff.t8 85.1574
R5027 start_buffer_0.start_buff.n9 start_buffer_0.start_buff.t5 83.8097
R5028 start_buffer_0.start_buff.n7 start_buffer_0.start_buff.t9 83.8097
R5029 start_buffer_0.start_buff.n18 start_buffer_0.start_buff.t2 83.7172
R5030 start_buffer_0.start_buff.n17 start_buffer_0.start_buff.t3 83.7172
R5031 start_buffer_0.start_buff.n20 start_buffer_0.start_buff.t1 83.7172
R5032 start_buffer_0.start_buff.n16 start_buffer_0.start_buff.t0 83.7172
R5033 start_buffer_0.start_buff.n5 start_buffer_0.start_buff.n3 36.1505
R5034 start_buffer_0.start_buff.n2 start_buffer_0.start_buff.n1 36.1505
R5035 start_buffer_0.start_buff.n5 start_buffer_0.start_buff.n4 34.5438
R5036 start_buffer_0.start_buff.n2 start_buffer_0.start_buff.n0 34.5438
R5037 start_buffer_0.start_buff.n8 start_buffer_0.start_buff.n6 11.8364
R5038 start_buffer_0.start_buff.n9 start_buffer_0.start_buff 8.40722
R5039 start_buffer_0.start_buff.n8 start_buffer_0.start_buff.n7 5.74235
R5040 start_buffer_0.start_buff.n19 start_buffer_0.start_buff.n17 5.16238
R5041 start_buffer_0.start_buff.n14 start_buffer_0.start_buff.n13 5.08518
R5042 start_buffer_0.start_buff start_buffer_0.start_buff.n16 4.70702
R5043 start_buffer_0.start_buff.n21 start_buffer_0.start_buff.n20 4.64452
R5044 start_buffer_0.start_buff.n19 start_buffer_0.start_buff.n18 4.64452
R5045 start_buffer_0.start_buff.n15 start_buffer_0.start_buff.n9 0.918978
R5046 start_buffer_0.start_buff.n21 start_buffer_0.start_buff.n19 0.518357
R5047 start_buffer_0.start_buff start_buffer_0.start_buff.n21 0.455857
R5048 start_buffer_0.start_buff.n16 start_buffer_0.start_buff.n15 0.3755
R5049 start_buffer_0.start_buff start_buffer_0.start_buff.n8 0.285656
R5050 start_buffer_0.start_buff.n15 start_buffer_0.start_buff.n14 0.247513
R5051 start_buffer_0.start_delay.n9 start_buffer_0.start_delay.t11 539.841
R5052 start_buffer_0.start_delay.n10 start_buffer_0.start_delay.t14 539.841
R5053 start_buffer_0.start_delay.n6 start_buffer_0.start_delay.t8 539.841
R5054 start_buffer_0.start_delay.n7 start_buffer_0.start_delay.t12 539.841
R5055 start_buffer_0.start_delay.n9 start_buffer_0.start_delay.t13 215.293
R5056 start_buffer_0.start_delay.n10 start_buffer_0.start_delay.t9 215.293
R5057 start_buffer_0.start_delay.n6 start_buffer_0.start_delay.t10 215.293
R5058 start_buffer_0.start_delay.n7 start_buffer_0.start_delay.t15 215.293
R5059 start_buffer_0.start_delay.n12 start_buffer_0.start_delay.n8 166.144
R5060 start_buffer_0.start_delay.n12 start_buffer_0.start_delay.n11 165.8
R5061 start_buffer_0.start_delay.n0 start_buffer_0.start_delay.t6 85.2499
R5062 start_buffer_0.start_delay.n1 start_buffer_0.start_delay.t5 85.2499
R5063 start_buffer_0.start_delay.n13 start_buffer_0.start_delay.t7 85.2499
R5064 start_buffer_0.start_delay.n3 start_buffer_0.start_delay.t4 84.7281
R5065 start_buffer_0.start_delay.n13 start_buffer_0.start_delay.t3 83.7172
R5066 start_buffer_0.start_delay.n0 start_buffer_0.start_delay.t2 83.7172
R5067 start_buffer_0.start_delay.n1 start_buffer_0.start_delay.t1 83.7172
R5068 start_buffer_0.start_delay.n4 start_buffer_0.start_delay.t0 83.7172
R5069 start_buffer_0.start_delay.n11 start_buffer_0.start_delay.n9 36.1505
R5070 start_buffer_0.start_delay.n8 start_buffer_0.start_delay.n6 36.1505
R5071 start_buffer_0.start_delay.n11 start_buffer_0.start_delay.n10 34.5438
R5072 start_buffer_0.start_delay.n8 start_buffer_0.start_delay.n7 34.5438
R5073 start_buffer_0.start_delay start_buffer_0.start_delay.n13 6.45821
R5074 start_buffer_0.start_delay.n2 start_buffer_0.start_delay.n0 5.16238
R5075 start_buffer_0.start_delay.n2 start_buffer_0.start_delay.n1 4.64452
R5076 start_buffer_0.start_delay.n5 start_buffer_0.start_delay.n4 4.64452
R5077 start_buffer_0.start_delay start_buffer_0.start_delay.n5 0.759429
R5078 start_buffer_0.start_delay start_buffer_0.start_delay.n12 0.53175
R5079 start_buffer_0.start_delay.n5 start_buffer_0.start_delay.n2 0.518357
R5080 start_buffer_0.start_delay.n4 start_buffer_0.start_delay.n3 0.3755
R5081 start_buffer_0.start_delay.n3 start_buffer_0.start_delay 0.234296
R5082 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 784.053
R5083 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 784.053
R5084 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 784.053
R5085 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 784.053
R5086 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 539.841
R5087 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 539.841
R5088 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 539.841
R5089 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 539.841
R5090 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 215.293
R5091 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 215.293
R5092 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 215.293
R5093 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 215.293
R5094 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 168.659
R5095 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 167.992
R5096 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 166.144
R5097 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 165.8
R5098 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 85.2499
R5099 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 85.2499
R5100 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 83.7172
R5101 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 83.7172
R5102 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 75.7282
R5103 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 66.3172
R5104 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 36.1505
R5105 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 36.1505
R5106 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 34.5438
R5107 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 34.5438
R5108 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 17.4005
R5109 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 17.4005
R5110 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 17.1141
R5111 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 9.52217
R5112 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 9.52217
R5113 vernier_delay_line_0.delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 6.45821
R5114 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 5.30824
R5115 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n15 4.94887
R5116 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 1.54347
R5117 vernier_delay_line_0.delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 1.06691
R5118 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 vernier_delay_line_0.delay_unit_2_0.in_2 0.602062
R5119 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd 0.453625
R5120 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n16 0.160656
R5121 a_n6458_3464.n28 a_n6458_3464.t13 543.053
R5122 a_n6458_3464.n26 a_n6458_3464.t21 543.053
R5123 a_n6458_3464.n24 a_n6458_3464.t32 543.053
R5124 a_n6458_3464.n22 a_n6458_3464.t10 543.053
R5125 a_n6458_3464.n20 a_n6458_3464.t17 543.053
R5126 a_n6458_3464.n18 a_n6458_3464.t30 543.053
R5127 a_n6458_3464.n16 a_n6458_3464.t8 543.053
R5128 a_n6458_3464.n14 a_n6458_3464.t19 543.053
R5129 a_n6458_3464.n12 a_n6458_3464.t26 543.053
R5130 a_n6458_3464.n10 a_n6458_3464.t37 543.053
R5131 a_n6458_3464.n8 a_n6458_3464.t15 543.053
R5132 a_n6458_3464.n6 a_n6458_3464.t23 543.053
R5133 a_n6458_3464.n4 a_n6458_3464.t33 543.053
R5134 a_n6458_3464.n2 a_n6458_3464.t11 543.053
R5135 a_n6458_3464.n1 a_n6458_3464.t28 543.053
R5136 a_n6458_3464.n0 a_n6458_3464.t35 543.053
R5137 a_n6458_3464.n28 a_n6458_3464.t16 221.72
R5138 a_n6458_3464.n26 a_n6458_3464.t24 221.72
R5139 a_n6458_3464.n24 a_n6458_3464.t34 221.72
R5140 a_n6458_3464.n22 a_n6458_3464.t12 221.72
R5141 a_n6458_3464.n20 a_n6458_3464.t20 221.72
R5142 a_n6458_3464.n18 a_n6458_3464.t31 221.72
R5143 a_n6458_3464.n16 a_n6458_3464.t9 221.72
R5144 a_n6458_3464.n14 a_n6458_3464.t22 221.72
R5145 a_n6458_3464.n12 a_n6458_3464.t27 221.72
R5146 a_n6458_3464.n10 a_n6458_3464.t39 221.72
R5147 a_n6458_3464.n8 a_n6458_3464.t18 221.72
R5148 a_n6458_3464.n6 a_n6458_3464.t25 221.72
R5149 a_n6458_3464.n4 a_n6458_3464.t36 221.72
R5150 a_n6458_3464.n2 a_n6458_3464.t14 221.72
R5151 a_n6458_3464.n1 a_n6458_3464.t29 221.72
R5152 a_n6458_3464.n0 a_n6458_3464.t38 221.72
R5153 a_n6458_3464.n3 a_n6458_3464.n1 218.32
R5154 a_n6458_3464.n29 a_n6458_3464.n28 217.734
R5155 a_n6458_3464.n27 a_n6458_3464.n26 217.734
R5156 a_n6458_3464.n25 a_n6458_3464.n24 217.734
R5157 a_n6458_3464.n23 a_n6458_3464.n22 217.734
R5158 a_n6458_3464.n21 a_n6458_3464.n20 217.734
R5159 a_n6458_3464.n19 a_n6458_3464.n18 217.734
R5160 a_n6458_3464.n17 a_n6458_3464.n16 217.734
R5161 a_n6458_3464.n15 a_n6458_3464.n14 217.734
R5162 a_n6458_3464.n13 a_n6458_3464.n12 217.734
R5163 a_n6458_3464.n11 a_n6458_3464.n10 217.734
R5164 a_n6458_3464.n9 a_n6458_3464.n8 217.734
R5165 a_n6458_3464.n7 a_n6458_3464.n6 217.734
R5166 a_n6458_3464.n5 a_n6458_3464.n4 217.734
R5167 a_n6458_3464.n3 a_n6458_3464.n2 217.734
R5168 a_n6458_3464.n30 a_n6458_3464.n0 213.234
R5169 a_n6458_3464.n35 a_n6458_3464.t5 85.2499
R5170 a_n6458_3464.n33 a_n6458_3464.t4 85.2499
R5171 a_n6458_3464.t7 a_n6458_3464.n37 85.2499
R5172 a_n6458_3464.n31 a_n6458_3464.t6 84.7173
R5173 a_n6458_3464.n37 a_n6458_3464.t2 83.7172
R5174 a_n6458_3464.n35 a_n6458_3464.t0 83.7172
R5175 a_n6458_3464.n33 a_n6458_3464.t3 83.7172
R5176 a_n6458_3464.n32 a_n6458_3464.t1 83.7172
R5177 a_n6458_3464.n36 a_n6458_3464.n35 5.16238
R5178 a_n6458_3464.n34 a_n6458_3464.n32 5.16238
R5179 a_n6458_3464.n30 a_n6458_3464.n29 5.08518
R5180 a_n6458_3464.n34 a_n6458_3464.n33 4.64452
R5181 a_n6458_3464.n37 a_n6458_3464.n36 4.64452
R5182 a_n6458_3464.n5 a_n6458_3464.n3 0.585177
R5183 a_n6458_3464.n7 a_n6458_3464.n5 0.585177
R5184 a_n6458_3464.n9 a_n6458_3464.n7 0.585177
R5185 a_n6458_3464.n11 a_n6458_3464.n9 0.585177
R5186 a_n6458_3464.n13 a_n6458_3464.n11 0.585177
R5187 a_n6458_3464.n15 a_n6458_3464.n13 0.585177
R5188 a_n6458_3464.n17 a_n6458_3464.n15 0.585177
R5189 a_n6458_3464.n19 a_n6458_3464.n17 0.585177
R5190 a_n6458_3464.n21 a_n6458_3464.n19 0.585177
R5191 a_n6458_3464.n23 a_n6458_3464.n21 0.585177
R5192 a_n6458_3464.n25 a_n6458_3464.n23 0.585177
R5193 a_n6458_3464.n27 a_n6458_3464.n25 0.585177
R5194 a_n6458_3464.n29 a_n6458_3464.n27 0.585177
R5195 a_n6458_3464.n36 a_n6458_3464.n34 0.518357
R5196 a_n6458_3464.n32 a_n6458_3464.n31 0.36463
R5197 a_n6458_3464.n31 a_n6458_3464.n30 0.226306
R5198 diff_gen_0.delay_unit_2_1.in_2.n3 diff_gen_0.delay_unit_2_1.in_2.t11 539.841
R5199 diff_gen_0.delay_unit_2_1.in_2.n4 diff_gen_0.delay_unit_2_1.in_2.t14 539.841
R5200 diff_gen_0.delay_unit_2_1.in_2.n0 diff_gen_0.delay_unit_2_1.in_2.t10 539.841
R5201 diff_gen_0.delay_unit_2_1.in_2.n1 diff_gen_0.delay_unit_2_1.in_2.t15 539.841
R5202 diff_gen_0.delay_unit_2_1.in_2.n3 diff_gen_0.delay_unit_2_1.in_2.t13 215.293
R5203 diff_gen_0.delay_unit_2_1.in_2.n4 diff_gen_0.delay_unit_2_1.in_2.t8 215.293
R5204 diff_gen_0.delay_unit_2_1.in_2.n0 diff_gen_0.delay_unit_2_1.in_2.t12 215.293
R5205 diff_gen_0.delay_unit_2_1.in_2.n1 diff_gen_0.delay_unit_2_1.in_2.t9 215.293
R5206 diff_gen_0.delay_unit_2_1.in_2.n6 diff_gen_0.delay_unit_2_1.in_2.n2 166.144
R5207 diff_gen_0.delay_unit_2_1.in_2.n6 diff_gen_0.delay_unit_2_1.in_2.n5 165.8
R5208 diff_gen_0.delay_unit_2_1.in_2.n7 diff_gen_0.delay_unit_2_1.in_2.t7 85.2499
R5209 diff_gen_0.delay_unit_2_1.in_2.n12 diff_gen_0.delay_unit_2_1.in_2.t6 85.2499
R5210 diff_gen_0.delay_unit_2_1.in_2.n12 diff_gen_0.delay_unit_2_1.in_2.t2 83.7172
R5211 diff_gen_0.delay_unit_2_1.in_2.n7 diff_gen_0.delay_unit_2_1.in_2.t0 83.7172
R5212 diff_gen_0.delay_unit_2_1.in_2.n11 diff_gen_0.delay_unit_2_1.in_2.n9 75.7282
R5213 diff_gen_0.delay_unit_2_1.in_2.n11 diff_gen_0.delay_unit_2_1.in_2.n10 66.3172
R5214 diff_gen_0.delay_unit_2_1.in_2.n5 diff_gen_0.delay_unit_2_1.in_2.n3 36.1505
R5215 diff_gen_0.delay_unit_2_1.in_2.n2 diff_gen_0.delay_unit_2_1.in_2.n0 36.1505
R5216 diff_gen_0.delay_unit_2_1.in_2.n5 diff_gen_0.delay_unit_2_1.in_2.n4 34.5438
R5217 diff_gen_0.delay_unit_2_1.in_2.n2 diff_gen_0.delay_unit_2_1.in_2.n1 34.5438
R5218 diff_gen_0.delay_unit_2_1.in_2.n10 diff_gen_0.delay_unit_2_1.in_2.t3 17.4005
R5219 diff_gen_0.delay_unit_2_1.in_2.n10 diff_gen_0.delay_unit_2_1.in_2.t1 17.4005
R5220 diff_gen_0.delay_unit_2_1.in_2.n9 diff_gen_0.delay_unit_2_1.in_2.t4 9.52217
R5221 diff_gen_0.delay_unit_2_1.in_2.n9 diff_gen_0.delay_unit_2_1.in_2.t5 9.52217
R5222 diff_gen_0.delay_unit_2_1.in_2.n8 diff_gen_0.delay_unit_2_1.in_2.n7 6.45821
R5223 diff_gen_0.delay_unit_2_1.in_2.n13 diff_gen_0.delay_unit_2_1.in_2.n11 5.30824
R5224 diff_gen_0.delay_unit_2_1.in_2.n13 diff_gen_0.delay_unit_2_1.in_2.n12 4.94887
R5225 diff_gen_0.delay_unit_2_1.in_2.n8 diff_gen_0.delay_unit_2_1.in_2.n6 1.06691
R5226 diff_gen_0.delay_unit_2_0.out_2 diff_gen_0.delay_unit_2_1.in_2.n8 0.188
R5227 diff_gen_0.delay_unit_2_0.out_2 diff_gen_0.delay_unit_2_1.in_2.n13 0.160656
R5228 diff_gen_0.delay_unit_2_1.in_1.n3 diff_gen_0.delay_unit_2_1.in_1.t11 539.841
R5229 diff_gen_0.delay_unit_2_1.in_1.n4 diff_gen_0.delay_unit_2_1.in_1.t9 539.841
R5230 diff_gen_0.delay_unit_2_1.in_1.n0 diff_gen_0.delay_unit_2_1.in_1.t10 539.841
R5231 diff_gen_0.delay_unit_2_1.in_1.n1 diff_gen_0.delay_unit_2_1.in_1.t15 539.841
R5232 diff_gen_0.delay_unit_2_1.in_1.n3 diff_gen_0.delay_unit_2_1.in_1.t14 215.293
R5233 diff_gen_0.delay_unit_2_1.in_1.n4 diff_gen_0.delay_unit_2_1.in_1.t12 215.293
R5234 diff_gen_0.delay_unit_2_1.in_1.n0 diff_gen_0.delay_unit_2_1.in_1.t13 215.293
R5235 diff_gen_0.delay_unit_2_1.in_1.n1 diff_gen_0.delay_unit_2_1.in_1.t8 215.293
R5236 diff_gen_0.delay_unit_2_1.in_1.n6 diff_gen_0.delay_unit_2_1.in_1.n2 166.149
R5237 diff_gen_0.delay_unit_2_1.in_1.n6 diff_gen_0.delay_unit_2_1.in_1.n5 165.8
R5238 diff_gen_0.delay_unit_2_1.in_1.n12 diff_gen_0.delay_unit_2_1.in_1.t4 85.1574
R5239 diff_gen_0.delay_unit_2_1.in_1.n7 diff_gen_0.delay_unit_2_1.in_1.t0 85.1574
R5240 diff_gen_0.delay_unit_2_1.in_1.n7 diff_gen_0.delay_unit_2_1.in_1.t1 83.8097
R5241 diff_gen_0.delay_unit_2_1.in_1.n12 diff_gen_0.delay_unit_2_1.in_1.t7 83.8097
R5242 diff_gen_0.delay_unit_2_1.in_1.n11 diff_gen_0.delay_unit_2_1.in_1.n10 74.288
R5243 diff_gen_0.delay_unit_2_1.in_1.n11 diff_gen_0.delay_unit_2_1.in_1.n9 67.7574
R5244 diff_gen_0.delay_unit_2_1.in_1.n5 diff_gen_0.delay_unit_2_1.in_1.n3 36.1505
R5245 diff_gen_0.delay_unit_2_1.in_1.n2 diff_gen_0.delay_unit_2_1.in_1.n1 36.1505
R5246 diff_gen_0.delay_unit_2_1.in_1.n5 diff_gen_0.delay_unit_2_1.in_1.n4 34.5438
R5247 diff_gen_0.delay_unit_2_1.in_1.n2 diff_gen_0.delay_unit_2_1.in_1.n0 34.5438
R5248 diff_gen_0.delay_unit_2_1.in_1.n9 diff_gen_0.delay_unit_2_1.in_1.t2 17.4005
R5249 diff_gen_0.delay_unit_2_1.in_1.n9 diff_gen_0.delay_unit_2_1.in_1.t3 17.4005
R5250 diff_gen_0.delay_unit_2_1.in_1.n8 diff_gen_0.delay_unit_2_1.in_1.n6 11.8364
R5251 diff_gen_0.delay_unit_2_1.in_1.n10 diff_gen_0.delay_unit_2_1.in_1.t5 9.52217
R5252 diff_gen_0.delay_unit_2_1.in_1.n10 diff_gen_0.delay_unit_2_1.in_1.t6 9.52217
R5253 diff_gen_0.delay_unit_2_1.in_1.n13 diff_gen_0.delay_unit_2_1.in_1.n11 5.83219
R5254 diff_gen_0.delay_unit_2_1.in_1.n8 diff_gen_0.delay_unit_2_1.in_1.n7 5.74235
R5255 diff_gen_0.delay_unit_2_1.in_1.n13 diff_gen_0.delay_unit_2_1.in_1.n12 5.49235
R5256 diff_gen_0.delay_unit_2_1.in_1 diff_gen_0.delay_unit_2_1.in_1.n13 1.32081
R5257 diff_gen_0.delay_unit_2_1.in_1 diff_gen_0.delay_unit_2_1.in_1.n8 0.285656
R5258 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 572.12
R5259 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 572.12
R5260 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 572.12
R5261 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 572.12
R5262 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 539.841
R5263 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 539.841
R5264 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 539.841
R5265 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 539.841
R5266 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 215.293
R5267 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 215.293
R5268 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 215.293
R5269 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 215.293
R5270 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 166.468
R5271 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 166.149
R5272 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 165.8
R5273 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 165.8
R5274 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 85.1574
R5275 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 83.8097
R5276 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 83.8097
R5277 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 83.7172
R5278 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 74.288
R5279 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 67.7574
R5280 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 36.1505
R5281 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 36.1505
R5282 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 34.5438
R5283 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 34.5438
R5284 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 17.4005
R5285 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 17.4005
R5286 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 16.0275
R5287 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 11.8364
R5288 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 9.52217
R5289 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 9.52217
R5290 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 6.02878
R5291 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 5.83219
R5292 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 5.74235
R5293 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 5.49235
R5294 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 1.44072
R5295 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 1.32081
R5296 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 784.053
R5297 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 784.053
R5298 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 784.053
R5299 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 784.053
R5300 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 539.841
R5301 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 539.841
R5302 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 539.841
R5303 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 539.841
R5304 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 215.293
R5305 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 215.293
R5306 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 215.293
R5307 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 215.293
R5308 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 168.659
R5309 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 167.992
R5310 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 166.144
R5311 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 165.8
R5312 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 85.2499
R5313 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 85.2499
R5314 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 83.7172
R5315 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 83.7172
R5316 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 75.7282
R5317 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 66.3172
R5318 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 36.1505
R5319 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 36.1505
R5320 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 34.5438
R5321 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 34.5438
R5322 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 17.4005
R5323 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 17.4005
R5324 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 17.1141
R5325 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 9.52217
R5326 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 9.52217
R5327 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 6.45821
R5328 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 5.30824
R5329 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 4.94887
R5330 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 1.70362
R5331 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 1.06691
R5332 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n15 0.602062
R5333 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.453625
R5334 diff_gen_0.delay_unit_2_4.in_1.n3 diff_gen_0.delay_unit_2_4.in_1.t14 539.841
R5335 diff_gen_0.delay_unit_2_4.in_1.n4 diff_gen_0.delay_unit_2_4.in_1.t10 539.841
R5336 diff_gen_0.delay_unit_2_4.in_1.n0 diff_gen_0.delay_unit_2_4.in_1.t13 539.841
R5337 diff_gen_0.delay_unit_2_4.in_1.n1 diff_gen_0.delay_unit_2_4.in_1.t9 539.841
R5338 diff_gen_0.delay_unit_2_4.in_1.n3 diff_gen_0.delay_unit_2_4.in_1.t8 215.293
R5339 diff_gen_0.delay_unit_2_4.in_1.n4 diff_gen_0.delay_unit_2_4.in_1.t12 215.293
R5340 diff_gen_0.delay_unit_2_4.in_1.n0 diff_gen_0.delay_unit_2_4.in_1.t15 215.293
R5341 diff_gen_0.delay_unit_2_4.in_1.n1 diff_gen_0.delay_unit_2_4.in_1.t11 215.293
R5342 diff_gen_0.delay_unit_2_4.in_1.n6 diff_gen_0.delay_unit_2_4.in_1.n2 166.149
R5343 diff_gen_0.delay_unit_2_4.in_1.n6 diff_gen_0.delay_unit_2_4.in_1.n5 165.8
R5344 diff_gen_0.delay_unit_2_4.in_1.n12 diff_gen_0.delay_unit_2_4.in_1.t2 85.1574
R5345 diff_gen_0.delay_unit_2_4.in_1.n7 diff_gen_0.delay_unit_2_4.in_1.t0 85.1574
R5346 diff_gen_0.delay_unit_2_4.in_1.n12 diff_gen_0.delay_unit_2_4.in_1.t5 83.8097
R5347 diff_gen_0.delay_unit_2_4.in_1.n7 diff_gen_0.delay_unit_2_4.in_1.t7 83.8097
R5348 diff_gen_0.delay_unit_2_4.in_1.n11 diff_gen_0.delay_unit_2_4.in_1.n10 74.288
R5349 diff_gen_0.delay_unit_2_4.in_1.n11 diff_gen_0.delay_unit_2_4.in_1.n9 67.7574
R5350 diff_gen_0.delay_unit_2_4.in_1.n5 diff_gen_0.delay_unit_2_4.in_1.n3 36.1505
R5351 diff_gen_0.delay_unit_2_4.in_1.n2 diff_gen_0.delay_unit_2_4.in_1.n1 36.1505
R5352 diff_gen_0.delay_unit_2_4.in_1.n5 diff_gen_0.delay_unit_2_4.in_1.n4 34.5438
R5353 diff_gen_0.delay_unit_2_4.in_1.n2 diff_gen_0.delay_unit_2_4.in_1.n0 34.5438
R5354 diff_gen_0.delay_unit_2_4.in_1.n9 diff_gen_0.delay_unit_2_4.in_1.t3 17.4005
R5355 diff_gen_0.delay_unit_2_4.in_1.n9 diff_gen_0.delay_unit_2_4.in_1.t1 17.4005
R5356 diff_gen_0.delay_unit_2_4.in_1.n8 diff_gen_0.delay_unit_2_4.in_1.n6 11.8364
R5357 diff_gen_0.delay_unit_2_4.in_1.n10 diff_gen_0.delay_unit_2_4.in_1.t6 9.52217
R5358 diff_gen_0.delay_unit_2_4.in_1.n10 diff_gen_0.delay_unit_2_4.in_1.t4 9.52217
R5359 diff_gen_0.delay_unit_2_4.in_1.n13 diff_gen_0.delay_unit_2_4.in_1.n11 5.83219
R5360 diff_gen_0.delay_unit_2_4.in_1.n8 diff_gen_0.delay_unit_2_4.in_1.n7 5.74235
R5361 diff_gen_0.delay_unit_2_4.in_1.n13 diff_gen_0.delay_unit_2_4.in_1.n12 5.49235
R5362 diff_gen_0.delay_unit_2_4.in_1 diff_gen_0.delay_unit_2_4.in_1.n13 1.32081
R5363 diff_gen_0.delay_unit_2_4.in_1 diff_gen_0.delay_unit_2_4.in_1.n8 0.285656
R5364 vernier_delay_line_0.start_neg.n3 vernier_delay_line_0.start_neg.t11 539.841
R5365 vernier_delay_line_0.start_neg.n4 vernier_delay_line_0.start_neg.t15 539.841
R5366 vernier_delay_line_0.start_neg.n0 vernier_delay_line_0.start_neg.t12 539.841
R5367 vernier_delay_line_0.start_neg.n1 vernier_delay_line_0.start_neg.t8 539.841
R5368 vernier_delay_line_0.start_neg.n3 vernier_delay_line_0.start_neg.t13 215.293
R5369 vernier_delay_line_0.start_neg.n4 vernier_delay_line_0.start_neg.t9 215.293
R5370 vernier_delay_line_0.start_neg.n0 vernier_delay_line_0.start_neg.t14 215.293
R5371 vernier_delay_line_0.start_neg.n1 vernier_delay_line_0.start_neg.t10 215.293
R5372 vernier_delay_line_0.start_neg.n6 vernier_delay_line_0.start_neg.n2 166.144
R5373 vernier_delay_line_0.start_neg.n6 vernier_delay_line_0.start_neg.n5 165.8
R5374 vernier_delay_line_0.start_neg.n11 vernier_delay_line_0.start_neg.t4 85.2499
R5375 vernier_delay_line_0.start_neg.n7 vernier_delay_line_0.start_neg.t6 85.2499
R5376 vernier_delay_line_0.start_neg.n11 vernier_delay_line_0.start_neg.t2 83.7172
R5377 vernier_delay_line_0.start_neg.n7 vernier_delay_line_0.start_neg.t7 83.7172
R5378 vernier_delay_line_0.start_neg.n10 vernier_delay_line_0.start_neg.n8 75.7282
R5379 vernier_delay_line_0.start_neg.n10 vernier_delay_line_0.start_neg.n9 66.3172
R5380 vernier_delay_line_0.start_neg.n5 vernier_delay_line_0.start_neg.n3 36.1505
R5381 vernier_delay_line_0.start_neg.n2 vernier_delay_line_0.start_neg.n0 36.1505
R5382 vernier_delay_line_0.start_neg.n5 vernier_delay_line_0.start_neg.n4 34.5438
R5383 vernier_delay_line_0.start_neg.n2 vernier_delay_line_0.start_neg.n1 34.5438
R5384 vernier_delay_line_0.start_neg.n9 vernier_delay_line_0.start_neg.t0 17.4005
R5385 vernier_delay_line_0.start_neg.n9 vernier_delay_line_0.start_neg.t1 17.4005
R5386 vernier_delay_line_0.start_neg.n8 vernier_delay_line_0.start_neg.t5 9.52217
R5387 vernier_delay_line_0.start_neg.n8 vernier_delay_line_0.start_neg.t3 9.52217
R5388 vernier_delay_line_0.start_neg vernier_delay_line_0.start_neg.n7 6.45821
R5389 vernier_delay_line_0.start_neg.n12 vernier_delay_line_0.start_neg.n10 5.30824
R5390 vernier_delay_line_0.start_neg.n12 vernier_delay_line_0.start_neg.n11 4.94887
R5391 vernier_delay_line_0.start_neg vernier_delay_line_0.start_neg.n6 0.754406
R5392 vernier_delay_line_0.start_neg vernier_delay_line_0.start_neg.n12 0.160656
R5393 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 784.053
R5394 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 784.053
R5395 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 784.053
R5396 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 784.053
R5397 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 539.841
R5398 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 539.841
R5399 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 539.841
R5400 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 539.841
R5401 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 215.293
R5402 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 215.293
R5403 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 215.293
R5404 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 215.293
R5405 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 168.659
R5406 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 167.992
R5407 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 166.144
R5408 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 165.8
R5409 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 85.2499
R5410 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 85.2499
R5411 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 83.7172
R5412 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 83.7172
R5413 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 75.7282
R5414 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 66.3172
R5415 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 36.1505
R5416 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 36.1505
R5417 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 34.5438
R5418 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 34.5438
R5419 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 17.4005
R5420 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 17.4005
R5421 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 17.1141
R5422 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 9.52217
R5423 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 9.52217
R5424 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 6.45821
R5425 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 5.30824
R5426 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 4.94887
R5427 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 1.70362
R5428 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 1.06691
R5429 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n15 0.602062
R5430 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.453625
R5431 a_5646_2192.n4 a_5646_2192.t12 32.0282
R5432 a_5646_2192.n9 a_5646_2192.n0 25.7663
R5433 a_5646_2192.n6 a_5646_2192.n1 25.75
R5434 a_5646_2192.n5 a_5646_2192.n2 25.75
R5435 a_5646_2192.n4 a_5646_2192.n3 25.75
R5436 a_5646_2192.n10 a_5646_2192.n9 25.288
R5437 a_5646_2192.n8 a_5646_2192.n7 24.288
R5438 a_5646_2192.n7 a_5646_2192.t2 5.8005
R5439 a_5646_2192.n7 a_5646_2192.t11 5.8005
R5440 a_5646_2192.n1 a_5646_2192.t10 5.8005
R5441 a_5646_2192.n1 a_5646_2192.t6 5.8005
R5442 a_5646_2192.n2 a_5646_2192.t7 5.8005
R5443 a_5646_2192.n2 a_5646_2192.t8 5.8005
R5444 a_5646_2192.n3 a_5646_2192.t9 5.8005
R5445 a_5646_2192.n3 a_5646_2192.t5 5.8005
R5446 a_5646_2192.n0 a_5646_2192.t0 5.8005
R5447 a_5646_2192.n0 a_5646_2192.t3 5.8005
R5448 a_5646_2192.n10 a_5646_2192.t1 5.8005
R5449 a_5646_2192.t4 a_5646_2192.n10 5.8005
R5450 a_5646_2192.n8 a_5646_2192.n6 1.94072
R5451 a_5646_2192.n9 a_5646_2192.n8 1.47876
R5452 a_5646_2192.n6 a_5646_2192.n5 0.478761
R5453 a_5646_2192.n5 a_5646_2192.n4 0.478761
R5454 a_5910_2192.n3 a_5910_2192.n2 34.9195
R5455 a_5910_2192.n2 a_5910_2192.n0 25.5407
R5456 a_5910_2192.n2 a_5910_2192.n1 25.2907
R5457 a_5910_2192.n0 a_5910_2192.t0 5.8005
R5458 a_5910_2192.n0 a_5910_2192.t1 5.8005
R5459 a_5910_2192.n1 a_5910_2192.t2 5.8005
R5460 a_5910_2192.n1 a_5910_2192.t3 5.8005
R5461 a_5910_2192.t4 a_5910_2192.n3 5.8005
R5462 a_5910_2192.n3 a_5910_2192.t5 5.8005
R5463 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 784.053
R5464 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 784.053
R5465 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 784.053
R5466 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 784.053
R5467 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 539.841
R5468 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 539.841
R5469 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 539.841
R5470 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 539.841
R5471 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 215.293
R5472 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 215.293
R5473 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 215.293
R5474 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 215.293
R5475 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 168.659
R5476 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 167.992
R5477 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 166.144
R5478 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 165.8
R5479 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 85.2499
R5480 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 85.2499
R5481 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 83.7172
R5482 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 83.7172
R5483 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 75.7282
R5484 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 66.3172
R5485 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 36.1505
R5486 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 36.1505
R5487 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 34.5438
R5488 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 34.5438
R5489 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 17.4005
R5490 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 17.4005
R5491 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 17.1141
R5492 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 9.52217
R5493 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 9.52217
R5494 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 6.45821
R5495 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 5.30824
R5496 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 4.94887
R5497 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 1.70362
R5498 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 1.06691
R5499 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 0.602062
R5500 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.453625
R5501 term_5.n1 term_5.t5 734.539
R5502 term_5.n1 term_5.t4 233.26
R5503 term_5.n2 term_5.n1 162.399
R5504 term_5.n2 term_5.n0 75.5108
R5505 term_5.n4 term_5.n3 66.3172
R5506 term_5.n3 term_5.t2 17.4005
R5507 term_5.n3 term_5.t0 17.4005
R5508 term_5.n0 term_5.t1 9.52217
R5509 term_5.n0 term_5.t3 9.52217
R5510 term_5 term_5.n4 5.08746
R5511 term_5.n4 term_5.n2 0.3755
R5512 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 572.12
R5513 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 572.12
R5514 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 572.12
R5515 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 572.12
R5516 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 539.841
R5517 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 539.841
R5518 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 539.841
R5519 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 539.841
R5520 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 215.293
R5521 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 215.293
R5522 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 215.293
R5523 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 215.293
R5524 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 166.468
R5525 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 166.149
R5526 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 165.8
R5527 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 165.8
R5528 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 85.1574
R5529 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 83.8097
R5530 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 83.8097
R5531 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 83.7172
R5532 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 74.288
R5533 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 67.7574
R5534 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 36.1505
R5535 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 36.1505
R5536 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 34.5438
R5537 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 34.5438
R5538 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 17.4005
R5539 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 17.4005
R5540 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 16.0275
R5541 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 11.8364
R5542 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 9.52217
R5543 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 9.52217
R5544 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 6.02878
R5545 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 5.83219
R5546 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 5.74235
R5547 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 5.49235
R5548 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 1.44072
R5549 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 1.32081
R5550 a_3364_2192.n4 a_3364_2192.t8 32.0282
R5551 a_3364_2192.n10 a_3364_2192.n9 25.7663
R5552 a_3364_2192.n6 a_3364_2192.n1 25.75
R5553 a_3364_2192.n5 a_3364_2192.n2 25.75
R5554 a_3364_2192.n4 a_3364_2192.n3 25.75
R5555 a_3364_2192.n9 a_3364_2192.n0 25.288
R5556 a_3364_2192.n8 a_3364_2192.n7 24.288
R5557 a_3364_2192.n7 a_3364_2192.t5 5.8005
R5558 a_3364_2192.n7 a_3364_2192.t11 5.8005
R5559 a_3364_2192.n1 a_3364_2192.t12 5.8005
R5560 a_3364_2192.n1 a_3364_2192.t9 5.8005
R5561 a_3364_2192.n2 a_3364_2192.t7 5.8005
R5562 a_3364_2192.n2 a_3364_2192.t1 5.8005
R5563 a_3364_2192.n3 a_3364_2192.t0 5.8005
R5564 a_3364_2192.n3 a_3364_2192.t10 5.8005
R5565 a_3364_2192.n0 a_3364_2192.t4 5.8005
R5566 a_3364_2192.n0 a_3364_2192.t2 5.8005
R5567 a_3364_2192.n10 a_3364_2192.t3 5.8005
R5568 a_3364_2192.t6 a_3364_2192.n10 5.8005
R5569 a_3364_2192.n8 a_3364_2192.n6 1.94072
R5570 a_3364_2192.n9 a_3364_2192.n8 1.47876
R5571 a_3364_2192.n6 a_3364_2192.n5 0.478761
R5572 a_3364_2192.n5 a_3364_2192.n4 0.478761
R5573 diff_gen_0.delay_unit_2_5.in_1.n3 diff_gen_0.delay_unit_2_5.in_1.t15 539.841
R5574 diff_gen_0.delay_unit_2_5.in_1.n4 diff_gen_0.delay_unit_2_5.in_1.t13 539.841
R5575 diff_gen_0.delay_unit_2_5.in_1.n0 diff_gen_0.delay_unit_2_5.in_1.t9 539.841
R5576 diff_gen_0.delay_unit_2_5.in_1.n1 diff_gen_0.delay_unit_2_5.in_1.t8 539.841
R5577 diff_gen_0.delay_unit_2_5.in_1.n3 diff_gen_0.delay_unit_2_5.in_1.t10 215.293
R5578 diff_gen_0.delay_unit_2_5.in_1.n4 diff_gen_0.delay_unit_2_5.in_1.t14 215.293
R5579 diff_gen_0.delay_unit_2_5.in_1.n0 diff_gen_0.delay_unit_2_5.in_1.t12 215.293
R5580 diff_gen_0.delay_unit_2_5.in_1.n1 diff_gen_0.delay_unit_2_5.in_1.t11 215.293
R5581 diff_gen_0.delay_unit_2_5.in_1.n6 diff_gen_0.delay_unit_2_5.in_1.n2 166.149
R5582 diff_gen_0.delay_unit_2_5.in_1.n6 diff_gen_0.delay_unit_2_5.in_1.n5 165.8
R5583 diff_gen_0.delay_unit_2_5.in_1.n12 diff_gen_0.delay_unit_2_5.in_1.t7 85.1574
R5584 diff_gen_0.delay_unit_2_5.in_1.n7 diff_gen_0.delay_unit_2_5.in_1.t3 85.1574
R5585 diff_gen_0.delay_unit_2_5.in_1.n12 diff_gen_0.delay_unit_2_5.in_1.t5 83.8097
R5586 diff_gen_0.delay_unit_2_5.in_1.n7 diff_gen_0.delay_unit_2_5.in_1.t4 83.8097
R5587 diff_gen_0.delay_unit_2_5.in_1.n11 diff_gen_0.delay_unit_2_5.in_1.n10 74.288
R5588 diff_gen_0.delay_unit_2_5.in_1.n11 diff_gen_0.delay_unit_2_5.in_1.n9 67.7574
R5589 diff_gen_0.delay_unit_2_5.in_1.n5 diff_gen_0.delay_unit_2_5.in_1.n3 36.1505
R5590 diff_gen_0.delay_unit_2_5.in_1.n2 diff_gen_0.delay_unit_2_5.in_1.n1 36.1505
R5591 diff_gen_0.delay_unit_2_5.in_1.n5 diff_gen_0.delay_unit_2_5.in_1.n4 34.5438
R5592 diff_gen_0.delay_unit_2_5.in_1.n2 diff_gen_0.delay_unit_2_5.in_1.n0 34.5438
R5593 diff_gen_0.delay_unit_2_5.in_1.n9 diff_gen_0.delay_unit_2_5.in_1.t2 17.4005
R5594 diff_gen_0.delay_unit_2_5.in_1.n9 diff_gen_0.delay_unit_2_5.in_1.t6 17.4005
R5595 diff_gen_0.delay_unit_2_5.in_1.n8 diff_gen_0.delay_unit_2_5.in_1.n6 11.8364
R5596 diff_gen_0.delay_unit_2_5.in_1.n10 diff_gen_0.delay_unit_2_5.in_1.t1 9.52217
R5597 diff_gen_0.delay_unit_2_5.in_1.n10 diff_gen_0.delay_unit_2_5.in_1.t0 9.52217
R5598 diff_gen_0.delay_unit_2_5.in_1.n13 diff_gen_0.delay_unit_2_5.in_1.n11 5.83219
R5599 diff_gen_0.delay_unit_2_5.in_1.n8 diff_gen_0.delay_unit_2_5.in_1.n7 5.74235
R5600 diff_gen_0.delay_unit_2_5.in_1.n13 diff_gen_0.delay_unit_2_5.in_1.n12 5.49235
R5601 diff_gen_0.delay_unit_2_4.out_1 diff_gen_0.delay_unit_2_5.in_1.n13 1.32081
R5602 diff_gen_0.delay_unit_2_4.out_1 diff_gen_0.delay_unit_2_5.in_1.n8 0.53175
R5603 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 879.481
R5604 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 742.783
R5605 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 665.16
R5606 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 623.388
R5607 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 523.774
R5608 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 431.807
R5609 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 427.875
R5610 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 357.26
R5611 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 208.537
R5612 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 168.077
R5613 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R5614 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 31.2347
R5615 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R5616 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 11.1806
R5617 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R5618 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 9.52217
R5619 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R5620 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R5621 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R5622 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 784.053
R5623 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 784.053
R5624 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 784.053
R5625 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 784.053
R5626 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 539.841
R5627 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 539.841
R5628 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 539.841
R5629 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 539.841
R5630 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 215.293
R5631 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 215.293
R5632 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 215.293
R5633 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 215.293
R5634 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 168.659
R5635 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 167.992
R5636 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 166.144
R5637 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 165.8
R5638 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 85.2499
R5639 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 85.2499
R5640 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 83.7172
R5641 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 83.7172
R5642 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 75.7282
R5643 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 66.3172
R5644 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 36.1505
R5645 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 36.1505
R5646 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 34.5438
R5647 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 34.5438
R5648 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 17.4005
R5649 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 17.4005
R5650 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 17.1141
R5651 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 9.52217
R5652 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 9.52217
R5653 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 6.45821
R5654 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 5.30824
R5655 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 4.94887
R5656 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 1.54347
R5657 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 1.06691
R5658 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n16 0.602062
R5659 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.453625
R5660 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n15 0.160656
R5661 a_15038_2192.n2 a_15038_2192.n1 34.9195
R5662 a_15038_2192.n2 a_15038_2192.n0 25.5407
R5663 a_15038_2192.n3 a_15038_2192.n2 25.2907
R5664 a_15038_2192.n1 a_15038_2192.t5 5.8005
R5665 a_15038_2192.n1 a_15038_2192.t3 5.8005
R5666 a_15038_2192.n0 a_15038_2192.t0 5.8005
R5667 a_15038_2192.n0 a_15038_2192.t1 5.8005
R5668 a_15038_2192.t4 a_15038_2192.n3 5.8005
R5669 a_15038_2192.n3 a_15038_2192.t2 5.8005
R5670 a_1082_2192.n4 a_1082_2192.t0 32.0282
R5671 a_1082_2192.n9 a_1082_2192.n0 25.7663
R5672 a_1082_2192.n6 a_1082_2192.n1 25.75
R5673 a_1082_2192.n5 a_1082_2192.n2 25.75
R5674 a_1082_2192.n4 a_1082_2192.n3 25.75
R5675 a_1082_2192.n10 a_1082_2192.n9 25.288
R5676 a_1082_2192.n8 a_1082_2192.n7 24.288
R5677 a_1082_2192.n7 a_1082_2192.t4 5.8005
R5678 a_1082_2192.n7 a_1082_2192.t2 5.8005
R5679 a_1082_2192.n1 a_1082_2192.t3 5.8005
R5680 a_1082_2192.n1 a_1082_2192.t12 5.8005
R5681 a_1082_2192.n2 a_1082_2192.t9 5.8005
R5682 a_1082_2192.n2 a_1082_2192.t11 5.8005
R5683 a_1082_2192.n3 a_1082_2192.t1 5.8005
R5684 a_1082_2192.n3 a_1082_2192.t10 5.8005
R5685 a_1082_2192.n0 a_1082_2192.t6 5.8005
R5686 a_1082_2192.n0 a_1082_2192.t5 5.8005
R5687 a_1082_2192.t8 a_1082_2192.n10 5.8005
R5688 a_1082_2192.n10 a_1082_2192.t7 5.8005
R5689 a_1082_2192.n8 a_1082_2192.n6 1.94072
R5690 a_1082_2192.n9 a_1082_2192.n8 1.47876
R5691 a_1082_2192.n6 a_1082_2192.n5 0.478761
R5692 a_1082_2192.n5 a_1082_2192.n4 0.478761
R5693 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 572.12
R5694 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 572.12
R5695 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 572.12
R5696 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 572.12
R5697 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 539.841
R5698 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 539.841
R5699 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 539.841
R5700 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 539.841
R5701 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 215.293
R5702 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 215.293
R5703 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 215.293
R5704 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 215.293
R5705 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 166.468
R5706 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 166.149
R5707 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 165.8
R5708 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 165.8
R5709 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 85.1574
R5710 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 83.8097
R5711 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 83.8097
R5712 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 83.7172
R5713 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 74.288
R5714 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 67.7574
R5715 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 36.1505
R5716 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 36.1505
R5717 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 34.5438
R5718 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 34.5438
R5719 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 17.4005
R5720 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 17.4005
R5721 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 16.0275
R5722 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 11.8364
R5723 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 9.52217
R5724 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 9.52217
R5725 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d 6.02878
R5726 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n17 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 5.83219
R5727 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 5.74235
R5728 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n17 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 5.49235
R5729 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 vernier_delay_line_0.delay_unit_2_0.in_1 2.20362
R5730 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 1.44072
R5731 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n17 1.32081
R5732 vernier_delay_line_0.delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 0.285656
R5733 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 572.12
R5734 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 572.12
R5735 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 572.12
R5736 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 572.12
R5737 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 539.841
R5738 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 539.841
R5739 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 539.841
R5740 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 539.841
R5741 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 215.293
R5742 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 215.293
R5743 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 215.293
R5744 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 215.293
R5745 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 166.468
R5746 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 166.149
R5747 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 165.8
R5748 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 165.8
R5749 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 85.1574
R5750 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 83.8097
R5751 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 83.8097
R5752 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 83.7172
R5753 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 74.288
R5754 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 67.7574
R5755 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 36.1505
R5756 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 36.1505
R5757 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 34.5438
R5758 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 34.5438
R5759 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 17.4005
R5760 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 17.4005
R5761 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 16.0275
R5762 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 11.8364
R5763 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 9.52217
R5764 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 9.52217
R5765 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 6.02878
R5766 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 5.83219
R5767 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 5.74235
R5768 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 5.49235
R5769 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 1.44072
R5770 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 1.32081
R5771 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 0.285656
R5772 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 784.053
R5773 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 784.053
R5774 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 784.053
R5775 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 784.053
R5776 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 539.841
R5777 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 539.841
R5778 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 539.841
R5779 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 539.841
R5780 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 215.293
R5781 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 215.293
R5782 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 215.293
R5783 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 215.293
R5784 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 168.659
R5785 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 167.992
R5786 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 166.144
R5787 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 165.8
R5788 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 85.2499
R5789 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 85.2499
R5790 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 83.7172
R5791 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 83.7172
R5792 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 75.7282
R5793 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 66.3172
R5794 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 36.1505
R5795 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 36.1505
R5796 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 34.5438
R5797 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 34.5438
R5798 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 17.4005
R5799 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 17.4005
R5800 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 17.1141
R5801 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 9.52217
R5802 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 9.52217
R5803 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 6.45821
R5804 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 5.30824
R5805 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 4.94887
R5806 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 1.70362
R5807 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 1.06691
R5808 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 0.602062
R5809 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.453625
R5810 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 890.727
R5811 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 742.783
R5812 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 665.16
R5813 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 623.388
R5814 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 523.774
R5815 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 431.807
R5816 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 427.875
R5817 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 364.733
R5818 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 208.5
R5819 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 168.007
R5820 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 75.2663
R5821 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 31.2728
R5822 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R5823 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R5824 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R5825 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 9.08234
R5826 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 8.00471
R5827 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 4.50239
R5828 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R5829 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 0.707022
R5830 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 879.481
R5831 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 742.783
R5832 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 665.16
R5833 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 623.388
R5834 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 523.774
R5835 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 431.807
R5836 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 427.875
R5837 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 357.26
R5838 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 208.537
R5839 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 168.077
R5840 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 75.5326
R5841 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R5842 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R5843 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 11.1806
R5844 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R5845 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R5846 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R5847 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R5848 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R5849 diff_gen_0.delay_unit_2_6.in_2.n3 diff_gen_0.delay_unit_2_6.in_2.t15 539.841
R5850 diff_gen_0.delay_unit_2_6.in_2.n4 diff_gen_0.delay_unit_2_6.in_2.t10 539.841
R5851 diff_gen_0.delay_unit_2_6.in_2.n0 diff_gen_0.delay_unit_2_6.in_2.t14 539.841
R5852 diff_gen_0.delay_unit_2_6.in_2.n1 diff_gen_0.delay_unit_2_6.in_2.t11 539.841
R5853 diff_gen_0.delay_unit_2_6.in_2.n3 diff_gen_0.delay_unit_2_6.in_2.t9 215.293
R5854 diff_gen_0.delay_unit_2_6.in_2.n4 diff_gen_0.delay_unit_2_6.in_2.t12 215.293
R5855 diff_gen_0.delay_unit_2_6.in_2.n0 diff_gen_0.delay_unit_2_6.in_2.t8 215.293
R5856 diff_gen_0.delay_unit_2_6.in_2.n1 diff_gen_0.delay_unit_2_6.in_2.t13 215.293
R5857 diff_gen_0.delay_unit_2_6.in_2.n6 diff_gen_0.delay_unit_2_6.in_2.n2 166.144
R5858 diff_gen_0.delay_unit_2_6.in_2.n6 diff_gen_0.delay_unit_2_6.in_2.n5 165.8
R5859 diff_gen_0.delay_unit_2_6.in_2.n12 diff_gen_0.delay_unit_2_6.in_2.t6 85.2499
R5860 diff_gen_0.delay_unit_2_6.in_2.n7 diff_gen_0.delay_unit_2_6.in_2.t1 85.2499
R5861 diff_gen_0.delay_unit_2_6.in_2.n12 diff_gen_0.delay_unit_2_6.in_2.t2 83.7172
R5862 diff_gen_0.delay_unit_2_6.in_2.n7 diff_gen_0.delay_unit_2_6.in_2.t0 83.7172
R5863 diff_gen_0.delay_unit_2_6.in_2.n11 diff_gen_0.delay_unit_2_6.in_2.n9 75.7282
R5864 diff_gen_0.delay_unit_2_6.in_2.n11 diff_gen_0.delay_unit_2_6.in_2.n10 66.3172
R5865 diff_gen_0.delay_unit_2_6.in_2.n5 diff_gen_0.delay_unit_2_6.in_2.n3 36.1505
R5866 diff_gen_0.delay_unit_2_6.in_2.n2 diff_gen_0.delay_unit_2_6.in_2.n0 36.1505
R5867 diff_gen_0.delay_unit_2_6.in_2.n5 diff_gen_0.delay_unit_2_6.in_2.n4 34.5438
R5868 diff_gen_0.delay_unit_2_6.in_2.n2 diff_gen_0.delay_unit_2_6.in_2.n1 34.5438
R5869 diff_gen_0.delay_unit_2_6.in_2.n10 diff_gen_0.delay_unit_2_6.in_2.t3 17.4005
R5870 diff_gen_0.delay_unit_2_6.in_2.n10 diff_gen_0.delay_unit_2_6.in_2.t4 17.4005
R5871 diff_gen_0.delay_unit_2_6.in_2.n9 diff_gen_0.delay_unit_2_6.in_2.t7 9.52217
R5872 diff_gen_0.delay_unit_2_6.in_2.n9 diff_gen_0.delay_unit_2_6.in_2.t5 9.52217
R5873 diff_gen_0.delay_unit_2_6.in_2.n8 diff_gen_0.delay_unit_2_6.in_2.n7 6.45821
R5874 diff_gen_0.delay_unit_2_6.in_2.n13 diff_gen_0.delay_unit_2_6.in_2.n11 5.30824
R5875 diff_gen_0.delay_unit_2_6.in_2.n13 diff_gen_0.delay_unit_2_6.in_2.n12 4.94887
R5876 diff_gen_0.delay_unit_2_6.in_2.n8 diff_gen_0.delay_unit_2_6.in_2.n6 1.06691
R5877 diff_gen_0.delay_unit_2_5.out_2 diff_gen_0.delay_unit_2_6.in_2.n8 0.188
R5878 diff_gen_0.delay_unit_2_5.out_2 diff_gen_0.delay_unit_2_6.in_2.n13 0.160656
R5879 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 572.12
R5880 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 572.12
R5881 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 572.12
R5882 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 572.12
R5883 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 539.841
R5884 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 539.841
R5885 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 539.841
R5886 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 539.841
R5887 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 215.293
R5888 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 215.293
R5889 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 215.293
R5890 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 215.293
R5891 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 166.468
R5892 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 166.149
R5893 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 165.8
R5894 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 165.8
R5895 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 85.1574
R5896 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 83.8097
R5897 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 83.8097
R5898 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 83.7172
R5899 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 74.288
R5900 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 67.7574
R5901 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 36.1505
R5902 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 36.1505
R5903 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 34.5438
R5904 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 34.5438
R5905 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 17.4005
R5906 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 17.4005
R5907 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 16.0275
R5908 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 11.8364
R5909 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 9.52217
R5910 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 9.52217
R5911 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 6.02878
R5912 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 5.83219
R5913 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 5.74235
R5914 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 5.49235
R5915 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 1.44072
R5916 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 1.32081
R5917 a_7928_2192.n4 a_7928_2192.t3 32.0282
R5918 a_7928_2192.n9 a_7928_2192.n0 25.7663
R5919 a_7928_2192.n6 a_7928_2192.n1 25.75
R5920 a_7928_2192.n5 a_7928_2192.n2 25.75
R5921 a_7928_2192.n4 a_7928_2192.n3 25.75
R5922 a_7928_2192.n10 a_7928_2192.n9 25.288
R5923 a_7928_2192.n8 a_7928_2192.n7 24.288
R5924 a_7928_2192.n7 a_7928_2192.t4 5.8005
R5925 a_7928_2192.n7 a_7928_2192.t9 5.8005
R5926 a_7928_2192.n1 a_7928_2192.t11 5.8005
R5927 a_7928_2192.n1 a_7928_2192.t0 5.8005
R5928 a_7928_2192.n2 a_7928_2192.t2 5.8005
R5929 a_7928_2192.n2 a_7928_2192.t12 5.8005
R5930 a_7928_2192.n3 a_7928_2192.t10 5.8005
R5931 a_7928_2192.n3 a_7928_2192.t1 5.8005
R5932 a_7928_2192.n0 a_7928_2192.t7 5.8005
R5933 a_7928_2192.n0 a_7928_2192.t6 5.8005
R5934 a_7928_2192.n10 a_7928_2192.t5 5.8005
R5935 a_7928_2192.t8 a_7928_2192.n10 5.8005
R5936 a_7928_2192.n8 a_7928_2192.n6 1.94072
R5937 a_7928_2192.n9 a_7928_2192.n8 1.47876
R5938 a_7928_2192.n6 a_7928_2192.n5 0.478761
R5939 a_7928_2192.n5 a_7928_2192.n4 0.478761
R5940 vernier_delay_line_0.start_pos.n3 vernier_delay_line_0.start_pos.t9 539.841
R5941 vernier_delay_line_0.start_pos.n4 vernier_delay_line_0.start_pos.t14 539.841
R5942 vernier_delay_line_0.start_pos.n0 vernier_delay_line_0.start_pos.t11 539.841
R5943 vernier_delay_line_0.start_pos.n1 vernier_delay_line_0.start_pos.t8 539.841
R5944 vernier_delay_line_0.start_pos.n3 vernier_delay_line_0.start_pos.t12 215.293
R5945 vernier_delay_line_0.start_pos.n4 vernier_delay_line_0.start_pos.t15 215.293
R5946 vernier_delay_line_0.start_pos.n0 vernier_delay_line_0.start_pos.t13 215.293
R5947 vernier_delay_line_0.start_pos.n1 vernier_delay_line_0.start_pos.t10 215.293
R5948 vernier_delay_line_0.start_pos.n6 vernier_delay_line_0.start_pos.n2 166.149
R5949 vernier_delay_line_0.start_pos.n6 vernier_delay_line_0.start_pos.n5 165.8
R5950 vernier_delay_line_0.start_pos.n12 vernier_delay_line_0.start_pos.t4 85.1574
R5951 vernier_delay_line_0.start_pos.n7 vernier_delay_line_0.start_pos.t0 85.1574
R5952 vernier_delay_line_0.start_pos.n12 vernier_delay_line_0.start_pos.t6 83.8097
R5953 vernier_delay_line_0.start_pos.n7 vernier_delay_line_0.start_pos.t1 83.8097
R5954 vernier_delay_line_0.start_pos.n11 vernier_delay_line_0.start_pos.n10 74.288
R5955 vernier_delay_line_0.start_pos.n11 vernier_delay_line_0.start_pos.n9 67.7574
R5956 vernier_delay_line_0.start_pos.n5 vernier_delay_line_0.start_pos.n3 36.1505
R5957 vernier_delay_line_0.start_pos.n2 vernier_delay_line_0.start_pos.n1 36.1505
R5958 vernier_delay_line_0.start_pos.n5 vernier_delay_line_0.start_pos.n4 34.5438
R5959 vernier_delay_line_0.start_pos.n2 vernier_delay_line_0.start_pos.n0 34.5438
R5960 vernier_delay_line_0.start_pos.n9 vernier_delay_line_0.start_pos.t2 17.4005
R5961 vernier_delay_line_0.start_pos.n9 vernier_delay_line_0.start_pos.t3 17.4005
R5962 vernier_delay_line_0.start_pos.n8 vernier_delay_line_0.start_pos.n6 11.8364
R5963 vernier_delay_line_0.start_pos.n10 vernier_delay_line_0.start_pos.t7 9.52217
R5964 vernier_delay_line_0.start_pos.n10 vernier_delay_line_0.start_pos.t5 9.52217
R5965 vernier_delay_line_0.start_pos.n13 vernier_delay_line_0.start_pos.n11 5.83219
R5966 vernier_delay_line_0.start_pos.n8 vernier_delay_line_0.start_pos.n7 5.74235
R5967 vernier_delay_line_0.start_pos.n13 vernier_delay_line_0.start_pos.n12 5.49235
R5968 vernier_delay_line_0.start_pos vernier_delay_line_0.start_pos.n13 1.32081
R5969 vernier_delay_line_0.start_pos vernier_delay_line_0.start_pos.n8 0.40675
R5970 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 784.053
R5971 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 784.053
R5972 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 784.053
R5973 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 784.053
R5974 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 539.841
R5975 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 539.841
R5976 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 539.841
R5977 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 539.841
R5978 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 215.293
R5979 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 215.293
R5980 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 215.293
R5981 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 215.293
R5982 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 168.659
R5983 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 167.992
R5984 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 166.144
R5985 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 165.8
R5986 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 85.2499
R5987 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 85.2499
R5988 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 83.7172
R5989 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 83.7172
R5990 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 75.7282
R5991 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 66.3172
R5992 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 36.1505
R5993 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 36.1505
R5994 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 34.5438
R5995 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 34.5438
R5996 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 17.4005
R5997 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 17.4005
R5998 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 17.1141
R5999 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 9.52217
R6000 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 9.52217
R6001 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 6.45821
R6002 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 5.30824
R6003 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 4.94887
R6004 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 1.54347
R6005 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 1.06691
R6006 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n16 0.602062
R6007 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.453625
R6008 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n15 0.160656
R6009 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 572.12
R6010 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 572.12
R6011 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 572.12
R6012 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 572.12
R6013 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 539.841
R6014 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 539.841
R6015 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 539.841
R6016 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 539.841
R6017 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 215.293
R6018 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 215.293
R6019 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 215.293
R6020 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 215.293
R6021 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 166.468
R6022 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 166.149
R6023 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 165.8
R6024 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 165.8
R6025 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 85.1574
R6026 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 83.8097
R6027 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 83.8097
R6028 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 83.7172
R6029 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 74.288
R6030 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 67.7574
R6031 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 36.1505
R6032 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 36.1505
R6033 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 34.5438
R6034 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 34.5438
R6035 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 17.4005
R6036 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 17.4005
R6037 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 16.0275
R6038 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 11.8364
R6039 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 9.52217
R6040 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 9.52217
R6041 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 6.02878
R6042 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 5.83219
R6043 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 5.74235
R6044 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 5.49235
R6045 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 1.44072
R6046 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 1.32081
R6047 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 0.285656
R6048 diff_gen_0.delay_unit_2_2.in_2.n3 diff_gen_0.delay_unit_2_2.in_2.t13 539.841
R6049 diff_gen_0.delay_unit_2_2.in_2.n4 diff_gen_0.delay_unit_2_2.in_2.t15 539.841
R6050 diff_gen_0.delay_unit_2_2.in_2.n0 diff_gen_0.delay_unit_2_2.in_2.t10 539.841
R6051 diff_gen_0.delay_unit_2_2.in_2.n1 diff_gen_0.delay_unit_2_2.in_2.t8 539.841
R6052 diff_gen_0.delay_unit_2_2.in_2.n3 diff_gen_0.delay_unit_2_2.in_2.t14 215.293
R6053 diff_gen_0.delay_unit_2_2.in_2.n4 diff_gen_0.delay_unit_2_2.in_2.t9 215.293
R6054 diff_gen_0.delay_unit_2_2.in_2.n0 diff_gen_0.delay_unit_2_2.in_2.t12 215.293
R6055 diff_gen_0.delay_unit_2_2.in_2.n1 diff_gen_0.delay_unit_2_2.in_2.t11 215.293
R6056 diff_gen_0.delay_unit_2_2.in_2.n6 diff_gen_0.delay_unit_2_2.in_2.n2 166.144
R6057 diff_gen_0.delay_unit_2_2.in_2.n6 diff_gen_0.delay_unit_2_2.in_2.n5 165.8
R6058 diff_gen_0.delay_unit_2_2.in_2.n7 diff_gen_0.delay_unit_2_2.in_2.t1 85.2499
R6059 diff_gen_0.delay_unit_2_2.in_2.n12 diff_gen_0.delay_unit_2_2.in_2.t7 85.2499
R6060 diff_gen_0.delay_unit_2_2.in_2.n12 diff_gen_0.delay_unit_2_2.in_2.t3 83.7172
R6061 diff_gen_0.delay_unit_2_2.in_2.n7 diff_gen_0.delay_unit_2_2.in_2.t0 83.7172
R6062 diff_gen_0.delay_unit_2_2.in_2.n11 diff_gen_0.delay_unit_2_2.in_2.n9 75.7282
R6063 diff_gen_0.delay_unit_2_2.in_2.n11 diff_gen_0.delay_unit_2_2.in_2.n10 66.3172
R6064 diff_gen_0.delay_unit_2_2.in_2.n5 diff_gen_0.delay_unit_2_2.in_2.n3 36.1505
R6065 diff_gen_0.delay_unit_2_2.in_2.n2 diff_gen_0.delay_unit_2_2.in_2.n0 36.1505
R6066 diff_gen_0.delay_unit_2_2.in_2.n5 diff_gen_0.delay_unit_2_2.in_2.n4 34.5438
R6067 diff_gen_0.delay_unit_2_2.in_2.n2 diff_gen_0.delay_unit_2_2.in_2.n1 34.5438
R6068 diff_gen_0.delay_unit_2_2.in_2.n10 diff_gen_0.delay_unit_2_2.in_2.t4 17.4005
R6069 diff_gen_0.delay_unit_2_2.in_2.n10 diff_gen_0.delay_unit_2_2.in_2.t2 17.4005
R6070 diff_gen_0.delay_unit_2_2.in_2.n9 diff_gen_0.delay_unit_2_2.in_2.t5 9.52217
R6071 diff_gen_0.delay_unit_2_2.in_2.n9 diff_gen_0.delay_unit_2_2.in_2.t6 9.52217
R6072 diff_gen_0.delay_unit_2_2.in_2.n8 diff_gen_0.delay_unit_2_2.in_2.n7 6.45821
R6073 diff_gen_0.delay_unit_2_2.in_2.n13 diff_gen_0.delay_unit_2_2.in_2.n11 5.30824
R6074 diff_gen_0.delay_unit_2_2.in_2.n13 diff_gen_0.delay_unit_2_2.in_2.n12 4.94887
R6075 diff_gen_0.delay_unit_2_2.in_2.n8 diff_gen_0.delay_unit_2_2.in_2.n6 1.06691
R6076 diff_gen_0.delay_unit_2_1.out_2 diff_gen_0.delay_unit_2_2.in_2.n8 0.188
R6077 diff_gen_0.delay_unit_2_1.out_2 diff_gen_0.delay_unit_2_2.in_2.n13 0.160656
R6078 diff_gen_0.delay_unit_2_3.in_1.n3 diff_gen_0.delay_unit_2_3.in_1.t12 539.841
R6079 diff_gen_0.delay_unit_2_3.in_1.n4 diff_gen_0.delay_unit_2_3.in_1.t8 539.841
R6080 diff_gen_0.delay_unit_2_3.in_1.n0 diff_gen_0.delay_unit_2_3.in_1.t11 539.841
R6081 diff_gen_0.delay_unit_2_3.in_1.n1 diff_gen_0.delay_unit_2_3.in_1.t15 539.841
R6082 diff_gen_0.delay_unit_2_3.in_1.n3 diff_gen_0.delay_unit_2_3.in_1.t14 215.293
R6083 diff_gen_0.delay_unit_2_3.in_1.n4 diff_gen_0.delay_unit_2_3.in_1.t10 215.293
R6084 diff_gen_0.delay_unit_2_3.in_1.n0 diff_gen_0.delay_unit_2_3.in_1.t13 215.293
R6085 diff_gen_0.delay_unit_2_3.in_1.n1 diff_gen_0.delay_unit_2_3.in_1.t9 215.293
R6086 diff_gen_0.delay_unit_2_3.in_1.n6 diff_gen_0.delay_unit_2_3.in_1.n2 166.149
R6087 diff_gen_0.delay_unit_2_3.in_1.n6 diff_gen_0.delay_unit_2_3.in_1.n5 165.8
R6088 diff_gen_0.delay_unit_2_3.in_1.n12 diff_gen_0.delay_unit_2_3.in_1.t1 85.1574
R6089 diff_gen_0.delay_unit_2_3.in_1.n7 diff_gen_0.delay_unit_2_3.in_1.t6 85.1574
R6090 diff_gen_0.delay_unit_2_3.in_1.n12 diff_gen_0.delay_unit_2_3.in_1.t4 83.8097
R6091 diff_gen_0.delay_unit_2_3.in_1.n7 diff_gen_0.delay_unit_2_3.in_1.t7 83.8097
R6092 diff_gen_0.delay_unit_2_3.in_1.n11 diff_gen_0.delay_unit_2_3.in_1.n10 74.288
R6093 diff_gen_0.delay_unit_2_3.in_1.n11 diff_gen_0.delay_unit_2_3.in_1.n9 67.7574
R6094 diff_gen_0.delay_unit_2_3.in_1.n5 diff_gen_0.delay_unit_2_3.in_1.n3 36.1505
R6095 diff_gen_0.delay_unit_2_3.in_1.n2 diff_gen_0.delay_unit_2_3.in_1.n1 36.1505
R6096 diff_gen_0.delay_unit_2_3.in_1.n5 diff_gen_0.delay_unit_2_3.in_1.n4 34.5438
R6097 diff_gen_0.delay_unit_2_3.in_1.n2 diff_gen_0.delay_unit_2_3.in_1.n0 34.5438
R6098 diff_gen_0.delay_unit_2_3.in_1.n9 diff_gen_0.delay_unit_2_3.in_1.t2 17.4005
R6099 diff_gen_0.delay_unit_2_3.in_1.n9 diff_gen_0.delay_unit_2_3.in_1.t0 17.4005
R6100 diff_gen_0.delay_unit_2_3.in_1.n8 diff_gen_0.delay_unit_2_3.in_1.n6 11.8364
R6101 diff_gen_0.delay_unit_2_3.in_1.n10 diff_gen_0.delay_unit_2_3.in_1.t5 9.52217
R6102 diff_gen_0.delay_unit_2_3.in_1.n10 diff_gen_0.delay_unit_2_3.in_1.t3 9.52217
R6103 diff_gen_0.delay_unit_2_3.in_1.n13 diff_gen_0.delay_unit_2_3.in_1.n11 5.83219
R6104 diff_gen_0.delay_unit_2_3.in_1.n8 diff_gen_0.delay_unit_2_3.in_1.n7 5.74235
R6105 diff_gen_0.delay_unit_2_3.in_1.n13 diff_gen_0.delay_unit_2_3.in_1.n12 5.49235
R6106 diff_gen_0.delay_unit_2_3.in_1 diff_gen_0.delay_unit_2_3.in_1.n13 1.32081
R6107 diff_gen_0.delay_unit_2_3.in_1 diff_gen_0.delay_unit_2_3.in_1.n8 0.285656
R6108 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 879.481
R6109 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 742.783
R6110 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 665.16
R6111 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 623.388
R6112 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 523.774
R6113 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 431.807
R6114 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 427.875
R6115 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 357.26
R6116 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 208.537
R6117 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 168.077
R6118 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 75.5326
R6119 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R6120 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R6121 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 11.1806
R6122 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 10.5958
R6123 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R6124 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R6125 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 0.803118
R6126 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 0.478761
R6127 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 572.12
R6128 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 572.12
R6129 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 572.12
R6130 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 572.12
R6131 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 539.841
R6132 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 539.841
R6133 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 539.841
R6134 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 539.841
R6135 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 215.293
R6136 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 215.293
R6137 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 215.293
R6138 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 215.293
R6139 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 166.468
R6140 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 166.149
R6141 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 165.8
R6142 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 165.8
R6143 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 85.1574
R6144 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 83.8097
R6145 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 83.8097
R6146 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 83.7172
R6147 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 74.288
R6148 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 67.7574
R6149 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 36.1505
R6150 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 36.1505
R6151 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 34.5438
R6152 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 34.5438
R6153 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 17.4005
R6154 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 17.4005
R6155 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 16.0275
R6156 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 11.8364
R6157 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 9.52217
R6158 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 9.52217
R6159 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 6.02878
R6160 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 5.83219
R6161 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 5.74235
R6162 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n17 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 5.49235
R6163 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 1.44072
R6164 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n17 1.32081
R6165 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 0.285656
R6166 a_17056_2192.n4 a_17056_2192.t1 32.0282
R6167 a_17056_2192.n9 a_17056_2192.n0 25.7663
R6168 a_17056_2192.n6 a_17056_2192.n1 25.75
R6169 a_17056_2192.n5 a_17056_2192.n2 25.75
R6170 a_17056_2192.n4 a_17056_2192.n3 25.75
R6171 a_17056_2192.n10 a_17056_2192.n9 25.288
R6172 a_17056_2192.n8 a_17056_2192.n7 24.288
R6173 a_17056_2192.n7 a_17056_2192.t8 5.8005
R6174 a_17056_2192.n7 a_17056_2192.t5 5.8005
R6175 a_17056_2192.n1 a_17056_2192.t4 5.8005
R6176 a_17056_2192.n1 a_17056_2192.t2 5.8005
R6177 a_17056_2192.n2 a_17056_2192.t0 5.8005
R6178 a_17056_2192.n2 a_17056_2192.t6 5.8005
R6179 a_17056_2192.n3 a_17056_2192.t7 5.8005
R6180 a_17056_2192.n3 a_17056_2192.t3 5.8005
R6181 a_17056_2192.n0 a_17056_2192.t9 5.8005
R6182 a_17056_2192.n0 a_17056_2192.t12 5.8005
R6183 a_17056_2192.t11 a_17056_2192.n10 5.8005
R6184 a_17056_2192.n10 a_17056_2192.t10 5.8005
R6185 a_17056_2192.n8 a_17056_2192.n6 1.94072
R6186 a_17056_2192.n9 a_17056_2192.n8 1.47876
R6187 a_17056_2192.n6 a_17056_2192.n5 0.478761
R6188 a_17056_2192.n5 a_17056_2192.n4 0.478761
R6189 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 890.727
R6190 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 742.783
R6191 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 665.16
R6192 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 623.388
R6193 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 523.774
R6194 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 431.807
R6195 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 427.875
R6196 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 364.733
R6197 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 208.5
R6198 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 168.007
R6199 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R6200 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 31.2728
R6201 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R6202 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R6203 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R6204 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 9.08234
R6205 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R6206 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R6207 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R6208 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R6209 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R6210 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 784.053
R6211 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 784.053
R6212 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 784.053
R6213 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 784.053
R6214 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 539.841
R6215 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 539.841
R6216 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 539.841
R6217 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 539.841
R6218 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 215.293
R6219 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 215.293
R6220 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 215.293
R6221 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 215.293
R6222 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 168.659
R6223 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 167.992
R6224 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 166.144
R6225 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 165.8
R6226 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 85.2499
R6227 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 85.2499
R6228 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 83.7172
R6229 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 83.7172
R6230 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 75.7282
R6231 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 66.3172
R6232 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 36.1505
R6233 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 36.1505
R6234 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 34.5438
R6235 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 34.5438
R6236 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 17.4005
R6237 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 17.4005
R6238 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 17.1141
R6239 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 9.52217
R6240 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 9.52217
R6241 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 6.45821
R6242 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 5.30824
R6243 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n15 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 4.94887
R6244 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 1.54347
R6245 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 1.06691
R6246 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n16 0.602062
R6247 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n16 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.453625
R6248 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n15 0.160656
R6249 a_10474_2192.n2 a_10474_2192.n1 34.9195
R6250 a_10474_2192.n3 a_10474_2192.n2 25.5407
R6251 a_10474_2192.n2 a_10474_2192.n0 25.2907
R6252 a_10474_2192.n1 a_10474_2192.t2 5.8005
R6253 a_10474_2192.n1 a_10474_2192.t1 5.8005
R6254 a_10474_2192.n0 a_10474_2192.t3 5.8005
R6255 a_10474_2192.n0 a_10474_2192.t0 5.8005
R6256 a_10474_2192.n3 a_10474_2192.t5 5.8005
R6257 a_10474_2192.t4 a_10474_2192.n3 5.8005
R6258 a_10210_2192.n4 a_10210_2192.t7 32.0282
R6259 a_10210_2192.n10 a_10210_2192.n9 25.7663
R6260 a_10210_2192.n6 a_10210_2192.n1 25.75
R6261 a_10210_2192.n5 a_10210_2192.n2 25.75
R6262 a_10210_2192.n4 a_10210_2192.n3 25.75
R6263 a_10210_2192.n9 a_10210_2192.n0 25.288
R6264 a_10210_2192.n8 a_10210_2192.n7 24.288
R6265 a_10210_2192.n7 a_10210_2192.t8 5.8005
R6266 a_10210_2192.n7 a_10210_2192.t2 5.8005
R6267 a_10210_2192.n1 a_10210_2192.t0 5.8005
R6268 a_10210_2192.n1 a_10210_2192.t4 5.8005
R6269 a_10210_2192.n2 a_10210_2192.t6 5.8005
R6270 a_10210_2192.n2 a_10210_2192.t3 5.8005
R6271 a_10210_2192.n3 a_10210_2192.t1 5.8005
R6272 a_10210_2192.n3 a_10210_2192.t5 5.8005
R6273 a_10210_2192.n0 a_10210_2192.t12 5.8005
R6274 a_10210_2192.n0 a_10210_2192.t9 5.8005
R6275 a_10210_2192.t11 a_10210_2192.n10 5.8005
R6276 a_10210_2192.n10 a_10210_2192.t10 5.8005
R6277 a_10210_2192.n8 a_10210_2192.n6 1.94072
R6278 a_10210_2192.n9 a_10210_2192.n8 1.47876
R6279 a_10210_2192.n6 a_10210_2192.n5 0.478761
R6280 a_10210_2192.n5 a_10210_2192.n4 0.478761
R6281 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 890.727
R6282 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 742.783
R6283 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 665.16
R6284 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 623.388
R6285 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 523.774
R6286 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 431.807
R6287 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 427.875
R6288 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 364.733
R6289 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 208.5
R6290 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 168.007
R6291 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R6292 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 31.2728
R6293 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 31.0337
R6294 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 9.52217
R6295 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R6296 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 9.08234
R6297 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R6298 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R6299 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R6300 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R6301 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R6302 a_8192_2192.n2 a_8192_2192.n1 34.9195
R6303 a_8192_2192.n2 a_8192_2192.n0 25.5407
R6304 a_8192_2192.n3 a_8192_2192.n2 25.2907
R6305 a_8192_2192.n1 a_8192_2192.t5 5.8005
R6306 a_8192_2192.n1 a_8192_2192.t3 5.8005
R6307 a_8192_2192.n0 a_8192_2192.t1 5.8005
R6308 a_8192_2192.n0 a_8192_2192.t0 5.8005
R6309 a_8192_2192.t4 a_8192_2192.n3 5.8005
R6310 a_8192_2192.n3 a_8192_2192.t2 5.8005
R6311 a_12756_2192.n3 a_12756_2192.n2 34.9195
R6312 a_12756_2192.n2 a_12756_2192.n0 25.5407
R6313 a_12756_2192.n2 a_12756_2192.n1 25.2907
R6314 a_12756_2192.n0 a_12756_2192.t4 5.8005
R6315 a_12756_2192.n0 a_12756_2192.t5 5.8005
R6316 a_12756_2192.n1 a_12756_2192.t0 5.8005
R6317 a_12756_2192.n1 a_12756_2192.t2 5.8005
R6318 a_12756_2192.t3 a_12756_2192.n3 5.8005
R6319 a_12756_2192.n3 a_12756_2192.t1 5.8005
R6320 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 890.727
R6321 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 742.783
R6322 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 665.16
R6323 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 623.388
R6324 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 523.774
R6325 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 431.807
R6326 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 427.875
R6327 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 364.733
R6328 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 208.5
R6329 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 168.007
R6330 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 75.2663
R6331 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 31.2728
R6332 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 31.0337
R6333 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R6334 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R6335 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 9.08234
R6336 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n8 8.00471
R6337 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n8 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 4.50239
R6338 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 0.898227
R6339 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 0.467891
R6340 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 0.23963
R6341 diff_gen_0.delay_unit_2_4.in_2.n3 diff_gen_0.delay_unit_2_4.in_2.t12 539.841
R6342 diff_gen_0.delay_unit_2_4.in_2.n4 diff_gen_0.delay_unit_2_4.in_2.t8 539.841
R6343 diff_gen_0.delay_unit_2_4.in_2.n0 diff_gen_0.delay_unit_2_4.in_2.t10 539.841
R6344 diff_gen_0.delay_unit_2_4.in_2.n1 diff_gen_0.delay_unit_2_4.in_2.t15 539.841
R6345 diff_gen_0.delay_unit_2_4.in_2.n3 diff_gen_0.delay_unit_2_4.in_2.t14 215.293
R6346 diff_gen_0.delay_unit_2_4.in_2.n4 diff_gen_0.delay_unit_2_4.in_2.t11 215.293
R6347 diff_gen_0.delay_unit_2_4.in_2.n0 diff_gen_0.delay_unit_2_4.in_2.t13 215.293
R6348 diff_gen_0.delay_unit_2_4.in_2.n1 diff_gen_0.delay_unit_2_4.in_2.t9 215.293
R6349 diff_gen_0.delay_unit_2_4.in_2.n6 diff_gen_0.delay_unit_2_4.in_2.n2 166.144
R6350 diff_gen_0.delay_unit_2_4.in_2.n6 diff_gen_0.delay_unit_2_4.in_2.n5 165.8
R6351 diff_gen_0.delay_unit_2_4.in_2.n7 diff_gen_0.delay_unit_2_4.in_2.t7 85.2499
R6352 diff_gen_0.delay_unit_2_4.in_2.n12 diff_gen_0.delay_unit_2_4.in_2.t5 85.2499
R6353 diff_gen_0.delay_unit_2_4.in_2.n12 diff_gen_0.delay_unit_2_4.in_2.t1 83.7172
R6354 diff_gen_0.delay_unit_2_4.in_2.n7 diff_gen_0.delay_unit_2_4.in_2.t6 83.7172
R6355 diff_gen_0.delay_unit_2_4.in_2.n11 diff_gen_0.delay_unit_2_4.in_2.n9 75.7282
R6356 diff_gen_0.delay_unit_2_4.in_2.n11 diff_gen_0.delay_unit_2_4.in_2.n10 66.3172
R6357 diff_gen_0.delay_unit_2_4.in_2.n5 diff_gen_0.delay_unit_2_4.in_2.n3 36.1505
R6358 diff_gen_0.delay_unit_2_4.in_2.n2 diff_gen_0.delay_unit_2_4.in_2.n0 36.1505
R6359 diff_gen_0.delay_unit_2_4.in_2.n5 diff_gen_0.delay_unit_2_4.in_2.n4 34.5438
R6360 diff_gen_0.delay_unit_2_4.in_2.n2 diff_gen_0.delay_unit_2_4.in_2.n1 34.5438
R6361 diff_gen_0.delay_unit_2_4.in_2.n10 diff_gen_0.delay_unit_2_4.in_2.t2 17.4005
R6362 diff_gen_0.delay_unit_2_4.in_2.n10 diff_gen_0.delay_unit_2_4.in_2.t0 17.4005
R6363 diff_gen_0.delay_unit_2_4.in_2.n9 diff_gen_0.delay_unit_2_4.in_2.t3 9.52217
R6364 diff_gen_0.delay_unit_2_4.in_2.n9 diff_gen_0.delay_unit_2_4.in_2.t4 9.52217
R6365 diff_gen_0.delay_unit_2_4.in_2.n8 diff_gen_0.delay_unit_2_4.in_2.n7 6.45821
R6366 diff_gen_0.delay_unit_2_4.in_2.n13 diff_gen_0.delay_unit_2_4.in_2.n11 5.30824
R6367 diff_gen_0.delay_unit_2_4.in_2.n13 diff_gen_0.delay_unit_2_4.in_2.n12 4.94887
R6368 diff_gen_0.delay_unit_2_4.in_2.n8 diff_gen_0.delay_unit_2_4.in_2.n6 1.06691
R6369 diff_gen_0.delay_unit_2_3.out_2 diff_gen_0.delay_unit_2_4.in_2.n8 0.188
R6370 diff_gen_0.delay_unit_2_3.out_2 diff_gen_0.delay_unit_2_4.in_2.n13 0.160656
R6371 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 890.727
R6372 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 742.783
R6373 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 665.16
R6374 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 623.388
R6375 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 523.774
R6376 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 431.807
R6377 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 427.875
R6378 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 364.733
R6379 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 208.5
R6380 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 168.007
R6381 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 75.2663
R6382 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 31.2728
R6383 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 31.0337
R6384 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R6385 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R6386 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 9.08234
R6387 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R6388 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 4.50239
R6389 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 0.898227
R6390 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 0.707022
R6391 term_2.n1 term_2.t5 734.539
R6392 term_2.n1 term_2.t4 233.26
R6393 term_2.n2 term_2.n1 162.399
R6394 term_2.n2 term_2.n0 75.5108
R6395 term_2.n4 term_2.n3 66.3172
R6396 term_2.n3 term_2.t2 17.4005
R6397 term_2.n3 term_2.t0 17.4005
R6398 term_2.n0 term_2.t1 9.52217
R6399 term_2.n0 term_2.t3 9.52217
R6400 term_2 term_2.n4 5.08746
R6401 term_2.n4 term_2.n2 0.3755
R6402 vernier_delay_line_0.delay_unit_2_0.out_1.n3 vernier_delay_line_0.delay_unit_2_0.out_1.t0 85.1574
R6403 vernier_delay_line_0.delay_unit_2_0.out_1.n3 vernier_delay_line_0.delay_unit_2_0.out_1.t4 83.8097
R6404 vernier_delay_line_0.delay_unit_2_0.out_1.n2 vernier_delay_line_0.delay_unit_2_0.out_1.n1 74.288
R6405 vernier_delay_line_0.delay_unit_2_0.out_1.n2 vernier_delay_line_0.delay_unit_2_0.out_1.n0 67.7574
R6406 vernier_delay_line_0.delay_unit_2_0.out_1.n0 vernier_delay_line_0.delay_unit_2_0.out_1.t2 17.4005
R6407 vernier_delay_line_0.delay_unit_2_0.out_1.n0 vernier_delay_line_0.delay_unit_2_0.out_1.t1 17.4005
R6408 vernier_delay_line_0.delay_unit_2_0.out_1.n1 vernier_delay_line_0.delay_unit_2_0.out_1.t3 9.52217
R6409 vernier_delay_line_0.delay_unit_2_0.out_1.n1 vernier_delay_line_0.delay_unit_2_0.out_1.t5 9.52217
R6410 vernier_delay_line_0.delay_unit_2_0.out_1.n4 vernier_delay_line_0.delay_unit_2_0.out_1.n2 5.83219
R6411 vernier_delay_line_0.delay_unit_2_0.out_1.n4 vernier_delay_line_0.delay_unit_2_0.out_1.n3 5.49235
R6412 vernier_delay_line_0.delay_unit_2_0.out_1 vernier_delay_line_0.delay_unit_2_0.out_1.n4 1.32081
R6413 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 879.481
R6414 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 742.783
R6415 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 665.16
R6416 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 623.388
R6417 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 523.774
R6418 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 431.807
R6419 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 427.875
R6420 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 357.26
R6421 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 208.537
R6422 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 168.077
R6423 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 75.5326
R6424 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R6425 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 31.2347
R6426 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 11.1806
R6427 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 10.5958
R6428 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 9.52217
R6429 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R6430 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 0.803118
R6431 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 0.23963
R6432 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 0.23963
R6433 a_3628_2192.n3 a_3628_2192.n2 34.9195
R6434 a_3628_2192.n2 a_3628_2192.n0 25.5407
R6435 a_3628_2192.n2 a_3628_2192.n1 25.2907
R6436 a_3628_2192.n0 a_3628_2192.t5 5.8005
R6437 a_3628_2192.n0 a_3628_2192.t4 5.8005
R6438 a_3628_2192.n1 a_3628_2192.t2 5.8005
R6439 a_3628_2192.n1 a_3628_2192.t0 5.8005
R6440 a_3628_2192.t3 a_3628_2192.n3 5.8005
R6441 a_3628_2192.n3 a_3628_2192.t1 5.8005
R6442 a_1346_2192.n2 a_1346_2192.n1 34.9195
R6443 a_1346_2192.n2 a_1346_2192.n0 25.5407
R6444 a_1346_2192.n3 a_1346_2192.n2 25.2907
R6445 a_1346_2192.n1 a_1346_2192.t3 5.8005
R6446 a_1346_2192.n1 a_1346_2192.t5 5.8005
R6447 a_1346_2192.n0 a_1346_2192.t0 5.8005
R6448 a_1346_2192.n0 a_1346_2192.t1 5.8005
R6449 a_1346_2192.n3 a_1346_2192.t2 5.8005
R6450 a_1346_2192.t4 a_1346_2192.n3 5.8005
R6451 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 890.727
R6452 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 742.783
R6453 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 665.16
R6454 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 623.388
R6455 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 523.774
R6456 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 431.807
R6457 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 427.875
R6458 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 364.733
R6459 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 208.5
R6460 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 168.007
R6461 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 75.2663
R6462 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 31.2728
R6463 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 31.0337
R6464 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 9.52217
R6465 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 9.52217
R6466 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 9.08234
R6467 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 8.00471
R6468 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 4.50239
R6469 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 0.898227
R6470 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 0.707022
R6471 term_4.n1 term_4.t5 734.539
R6472 term_4.n1 term_4.t4 233.26
R6473 term_4.n2 term_4.n1 162.399
R6474 term_4.n2 term_4.n0 75.5108
R6475 term_4.n4 term_4.n3 66.3172
R6476 term_4.n3 term_4.t3 17.4005
R6477 term_4.n3 term_4.t0 17.4005
R6478 term_4.n0 term_4.t1 9.52217
R6479 term_4.n0 term_4.t2 9.52217
R6480 term_4 term_4.n4 5.08746
R6481 term_4.n4 term_4.n2 0.3755
R6482 a_17320_2192.n3 a_17320_2192.n2 34.9195
R6483 a_17320_2192.n2 a_17320_2192.n0 25.5407
R6484 a_17320_2192.n2 a_17320_2192.n1 25.2907
R6485 a_17320_2192.n0 a_17320_2192.t5 5.8005
R6486 a_17320_2192.n0 a_17320_2192.t4 5.8005
R6487 a_17320_2192.n1 a_17320_2192.t2 5.8005
R6488 a_17320_2192.n1 a_17320_2192.t0 5.8005
R6489 a_17320_2192.t3 a_17320_2192.n3 5.8005
R6490 a_17320_2192.n3 a_17320_2192.t1 5.8005
R6491 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 879.481
R6492 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 742.783
R6493 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 665.16
R6494 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 623.388
R6495 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 523.774
R6496 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 431.807
R6497 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 427.875
R6498 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 357.26
R6499 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 208.537
R6500 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 168.077
R6501 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 75.5326
R6502 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n7 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 31.2347
R6503 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 31.2347
R6504 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 11.1806
R6505 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n7 10.5958
R6506 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 9.52217
R6507 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 9.52217
R6508 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 0.803118
R6509 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n7 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 0.23963
R6510 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 0.23963
R6511 term_1.n1 term_1.t5 734.539
R6512 term_1.n1 term_1.t4 233.26
R6513 term_1.n2 term_1.n1 162.399
R6514 term_1.n2 term_1.n0 75.5108
R6515 term_1.n4 term_1.n3 66.3172
R6516 term_1.n3 term_1.t3 17.4005
R6517 term_1.n3 term_1.t0 17.4005
R6518 term_1.n0 term_1.t1 9.52217
R6519 term_1.n0 term_1.t2 9.52217
R6520 term_1 term_1.n4 5.08746
R6521 term_1.n4 term_1.n2 0.3755
R6522 term_3.n1 term_3.t5 734.539
R6523 term_3.n1 term_3.t4 233.26
R6524 term_3.n2 term_3.n1 162.399
R6525 term_3.n2 term_3.n0 75.5108
R6526 term_3.n4 term_3.n3 66.3172
R6527 term_3.n3 term_3.t0 17.4005
R6528 term_3.n3 term_3.t2 17.4005
R6529 term_3.n0 term_3.t3 9.52217
R6530 term_3.n0 term_3.t1 9.52217
R6531 term_3 term_3.n4 5.08746
R6532 term_3.n4 term_3.n2 0.3755
R6533 term_0.n1 term_0.t5 734.539
R6534 term_0.n1 term_0.t4 233.26
R6535 term_0.n2 term_0.n1 162.399
R6536 term_0.n2 term_0.n0 75.5108
R6537 term_0.n4 term_0.n3 66.3172
R6538 term_0.n3 term_0.t0 17.4005
R6539 term_0.n3 term_0.t2 17.4005
R6540 term_0.n0 term_0.t3 9.52217
R6541 term_0.n0 term_0.t1 9.52217
R6542 term_0 term_0.n4 5.08746
R6543 term_0.n4 term_0.n2 0.3755
R6544 term_6.n1 term_6.t5 734.539
R6545 term_6.n1 term_6.t4 233.26
R6546 term_6.n2 term_6.n1 162.399
R6547 term_6.n2 term_6.n0 75.5108
R6548 term_6.n4 term_6.n3 66.3172
R6549 term_6.n3 term_6.t0 17.4005
R6550 term_6.n3 term_6.t2 17.4005
R6551 term_6.n0 term_6.t3 9.52217
R6552 term_6.n0 term_6.t1 9.52217
R6553 term_6 term_6.n4 5.08746
R6554 term_6.n4 term_6.n2 0.3755
R6555 start.n0 start.t0 543.053
R6556 start.n0 start.t1 221.72
R6557 start start.n0 213.398
R6558 stop.n0 stop.t0 543.053
R6559 stop.n0 stop.t1 221.72
R6560 stop stop.n0 213.398
C0 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.28924f
C1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VDD 0.706518f
C2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.501329f
C3 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 1.99e-19
C4 a_15162_296# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.005542f
C5 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.953579f
C6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.006183f
C7 a_17176_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.15e-21
C8 term_6 a_14894_160# 0.098219f
C9 a_17176_160# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.196688f
C10 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.132512f
C11 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.003768f
C12 a_8048_160# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.01482f
C13 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_5734_2192# 0.007929f
C14 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.019931f
C15 a_4130_730# term_1 0.013457f
C16 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.003768f
C17 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 VDD 5.07265f
C18 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_4168_1376# 7.19e-22
C19 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.237663f
C20 term_0 a_1886_1376# 0.014823f
C21 VDD vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 2.57087f
C22 a_8732_1376# a_8694_296# 1.02e-19
C23 term_5 a_13258_296# 0.005542f
C24 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 1.24e-19
C25 a_12612_160# a_13296_1376# 0.005826f
C26 term_1 a_3484_160# 0.098219f
C27 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1202_160# 0.164402f
C28 a_10598_730# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.003664f
C29 VDD a_5766_160# 1.42789f
C30 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15540_730# 0.504416f
C31 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_4168_1376# 2.36e-21
C32 VDD vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 3.23813f
C33 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17822_730# 0.504416f
C34 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.231672f
C35 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_4130_730# 0.033952f
C36 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.752988f
C37 a_10330_160# term_4 0.098219f
C38 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.59e-20
C39 vernier_delay_line_0.delay_unit_2_0.out_2 vernier_delay_line_0.delay_unit_2_0.out_1 0.031607f
C40 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_1886_1376# 0.162625f
C41 a_n8488_3464# a_n6748_3464# 5.08e-20
C42 VDD vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 2.43248f
C43 VDD a_n8198_3464# 1.1544f
C44 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_3484_160# 0.164402f
C45 a_6412_296# term_2 0.005542f
C46 VDD diff_gen_0.delay_unit_2_4.in_1 4.44104f
C47 a_3452_2192# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.09966f
C48 a_8048_160# VDD 1.42789f
C49 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_6034_730# 0.003664f
C50 VDD vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.706518f
C51 VDD vernier_delay_line_0.start_pos 4.75638f
C52 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 4.73e-19
C53 a_8316_730# term_3 0.492009f
C54 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.871529f
C55 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.006183f
C56 a_14862_2192# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.192064f
C57 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12880_296# 0.005542f
C58 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.001059f
C59 a_15540_296# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.174293f
C60 term_6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.201251f
C61 a_1470_296# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.005542f
C62 term_7 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.53e-22
C63 a_11014_1376# a_12612_160# 0.005973f
C64 VDD term_0 0.587468f
C65 a_17176_160# a_17144_2192# 2.08e-21
C66 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 1.17e-19
C67 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1848_730# 0.504416f
C68 term_7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.201251f
C69 a_12880_730# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.003664f
C70 VDD vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.57087f
C71 a_3752_296# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.005542f
C72 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 4.73e-19
C73 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.953579f
C74 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.747722f
C75 a_8732_1376# a_8694_730# 0.030083f
C76 term_6 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.53e-22
C77 term_4 a_11014_1376# 0.014823f
C78 VDD vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 2.57483f
C79 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.019931f
C80 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_12880_730# 0.013457f
C81 a_1170_2192# vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.007929f
C82 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_8016_2192# 0.192064f
C83 VDD diff_gen_0.delay_unit_2_3.in_1 4.44078f
C84 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17444_296# 0.005542f
C85 VDD vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.706518f
C86 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.59e-20
C87 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_4168_1376# 5.04e-20
C88 VDD diff_gen_0.delay_unit_2_6.in_1 4.42926f
C89 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.231672f
C90 a_n7908_3464# a_n6748_3464# 2.78e-19
C91 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 4.73e-19
C92 VDD vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 3.23801f
C93 a_13258_296# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.012202f
C94 VDD a_n7618_3464# 1.1544f
C95 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 term_3 0.10528f
C96 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.231672f
C97 VDD vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.706518f
C98 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.010157f
C99 a_5766_160# a_6034_730# 0.030392f
C100 VDD a_15578_1376# 1.40782f
C101 a_10976_730# a_10976_296# 0.003413f
C102 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.99e-19
C103 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_1 6.28e-22
C104 VDD a_4168_1376# 1.40782f
C105 start_buffer_0.start_buff a_n8778_3464# 6.61e-19
C106 a_4130_296# term_1 0.005542f
C107 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13258_296# 0.174293f
C108 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.237663f
C109 a_8732_1376# term_4 6.12e-20
C110 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.019931f
C111 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.99e-19
C112 a_8048_160# a_8016_2192# 2.08e-21
C113 VDD a_1886_1376# 1.40782f
C114 a_8732_1376# vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 5.04e-20
C115 a_13258_730# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.003607f
C116 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.747722f
C117 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_3752_730# 0.035356f
C118 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_8316_730# 1.47e-19
C119 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VDD 0.706518f
C120 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.132512f
C121 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_4130_730# 0.504416f
C122 a_10330_160# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.45e-19
C123 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.99e-19
C124 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.003768f
C125 term_5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 1.13e-20
C126 a_6412_296# a_6450_1376# 1.02e-19
C127 a_4130_296# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.012202f
C128 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.237663f
C129 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_3484_160# 0.01482f
C130 a_1170_2192# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 1.06381f
C131 a_17444_730# VDD 0.497771f
C132 VDD vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 5.07265f
C133 a_15162_296# a_15162_730# 0.003413f
C134 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_3484_160# 6.08e-20
C135 term_7 a_17822_296# 0.005542f
C136 term_6 a_15578_1376# 0.014823f
C137 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 VDD 3.23801f
C138 a_12580_2192# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.007929f
C139 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 a_10976_296# 0.012202f
C140 a_8694_296# term_3 0.005542f
C141 a_17860_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.162625f
C142 a_8048_160# a_8316_730# 0.030392f
C143 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_6034_730# 0.035356f
C144 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10598_730# 0.013457f
C145 start_buffer_0.start_delay diff_gen_0.delay_unit_2_1.in_1 0.401491f
C146 a_n7328_3464# a_n6748_3464# 0.001101f
C147 diff_gen_0.delay_unit_2_1.in_1 a_n7328_3464# 6.02e-19
C148 term_4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 1.13e-20
C149 VDD a_n7038_3464# 1.1544f
C150 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.871529f
C151 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 term_2 3.69e-19
C152 VDD a_12880_296# 6.18e-19
C153 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.138536f
C154 term_5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.201251f
C155 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 6.79e-20
C156 a_15162_730# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.003664f
C157 a_11014_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.36e-21
C158 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.006183f
C159 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 0.953579f
C160 term_6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.13e-20
C161 a_14894_160# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 3.45e-19
C162 a_14894_160# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 4.55e-19
C163 a_6450_1376# term_2 0.014823f
C164 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 1.17e-19
C165 a_n8778_3464# stop 0.072972f
C166 a_12612_160# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 4.55e-19
C167 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_6034_730# 0.013457f
C168 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_5766_160# 1.15e-21
C169 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.138536f
C170 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 a_6450_1376# 7.19e-22
C171 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 VDD 5.07265f
C172 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.018644f
C173 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 4.73e-19
C174 a_10330_160# a_11014_1376# 0.005826f
C175 VDD a_12880_730# 0.497771f
C176 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 4.73e-19
C177 a_17822_730# VDD 0.497547f
C178 a_12880_730# a_12880_296# 0.003413f
C179 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 a_1470_730# 1.47e-19
C180 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_6450_1376# 2.36e-21
C181 a_8048_160# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.164402f
C182 a_13296_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 3.26e-19
C183 a_5734_2192# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.09966f
C184 a_1470_296# a_1470_730# 0.003413f
C185 VDD vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.57087f
C186 term_6 VDD 0.587468f
C187 a_15578_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 3.26e-19
C188 a_6034_296# a_5766_160# 1.02e-19
C189 a_8694_730# term_3 0.013457f
C190 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.138536f
C191 a_8732_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.162625f
C192 a_1848_296# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.174293f
C193 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 a_1202_160# 4.55e-19
C194 a_3752_296# a_3752_730# 0.003413f
C195 term_4 a_10976_730# 0.013457f
C196 a_14894_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.01482f
C197 a_17176_160# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.01482f
C198 a_3752_296# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.010872f
C199 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.747722f
C200 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10598_296# 0.005542f
C201 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_0 6.28e-22
C202 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.001059f
C203 VDD a_13258_296# 6.18e-19
C204 a_4130_296# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.174293f
C205 a_n11872_5654# start_buffer_0.start_delay 7.1e-20
C206 a_17444_730# a_17444_296# 0.003413f
C207 a_6412_730# a_6412_296# 0.003413f
C208 a_17860_1376# a_17822_296# 1.02e-19
C209 a_8732_1376# a_10330_160# 0.005973f
C210 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8316_730# 0.013457f
C211 VDD a_10598_730# 0.497771f
C212 a_15540_730# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.033952f
C213 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 6.79e-20
C214 a_8316_296# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.010872f
C215 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C216 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.237663f
C217 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.752988f
C218 a_12612_160# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.15e-21
C219 a_17444_730# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.003664f
C220 term_5 a_12612_160# 0.098219f
C221 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 7.03e-19
C222 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 6.79e-20
C223 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.747722f
C224 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 6.79e-20
C225 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1470_730# 0.003664f
C226 a_17176_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.45e-19
C227 VDD a_6034_730# 0.497771f
C228 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_5766_160# 3.84e-19
C229 term_0 a_1202_160# 0.098219f
C230 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 9.61e-20
C231 a_n8778_3464# a_n8488_3464# 0.083149f
C232 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 term_3 3.69e-19
C233 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 4.28924f
C234 a_4168_1376# term_1 0.014823f
C235 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_6450_1376# 5.04e-20
C236 a_6034_296# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.010872f
C237 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 9.61e-20
C238 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.010157f
C239 a_17444_296# VDD 6.18e-19
C240 term_4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.10528f
C241 a_5734_2192# a_5766_160# 2.08e-21
C242 a_15540_296# a_15540_730# 0.003413f
C243 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.018644f
C244 term_1 a_1886_1376# 6.12e-20
C245 a_15540_296# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.012202f
C246 VDD vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 2.43248f
C247 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.132512f
C248 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_1202_160# 0.196688f
C249 a_10598_730# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.035356f
C250 a_8316_730# VDD 0.497771f
C251 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.871529f
C252 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_4168_1376# 0.197073f
C253 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 9.61e-20
C254 a_10330_160# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 3.84e-19
C255 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.132512f
C256 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_4130_730# 0.003607f
C257 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.231672f
C258 term_7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq 0.229061f
C259 a_3752_730# a_3484_160# 0.030392f
C260 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_1886_1376# 3.26e-19
C261 a_6412_730# term_2 0.013457f
C262 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_5766_160# 6.08e-20
C263 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10976_296# 0.174293f
C264 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_3484_160# 0.196688f
C265 a_6034_296# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.005542f
C266 a_12580_2192# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.09966f
C267 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 term_1 3.69e-19
C268 a_3452_2192# vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 1.06381f
C269 a_14862_2192# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.007929f
C270 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 1.24e-19
C271 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.501329f
C272 start_buffer_0.start_buff VDD 7.20373f
C273 a_17822_730# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.033952f
C274 VDD a_10598_296# 6.18e-19
C275 term_6 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 6.28e-22
C276 a_6412_296# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.012202f
C277 a_1202_160# a_1886_1376# 0.005826f
C278 a_5734_2192# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 1.06381f
C279 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_17144_2192# 1.06381f
C280 VDD term_1 0.587468f
C281 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.441403f
C282 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.138536f
C283 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.006183f
C284 a_n8488_3464# a_n8198_3464# 0.083149f
C285 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.752988f
C286 a_10330_160# a_10298_2192# 2.08e-21
C287 VDD vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 2.43248f
C288 a_12612_160# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.164402f
C289 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.953579f
C290 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1848_730# 0.033952f
C291 a_15578_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.36e-21
C292 a_15578_1376# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 5.04e-20
C293 VDD vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 2.43248f
C294 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.001059f
C295 term_0 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.229061f
C296 a_13296_1376# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 5.04e-20
C297 a_13296_1376# a_13258_730# 0.030083f
C298 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8694_296# 0.174293f
C299 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 term_1 1.13e-20
C300 a_17176_160# a_15578_1376# 0.005973f
C301 a_12612_160# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.01482f
C302 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 a_10598_296# 0.010872f
C303 VDD vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 5.07265f
C304 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 2.59e-20
C305 term_4 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 6.28e-22
C306 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 term_3 0.201251f
C307 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.132512f
C308 a_6034_296# VDD 6.18e-19
C309 a_n11872_5654# start 0.076831f
C310 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.138536f
C311 VDD a_1202_160# 1.42748f
C312 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.747722f
C313 a_8048_160# vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 4.55e-19
C314 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 6.79e-20
C315 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_2 0.10528f
C316 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.010157f
C317 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.953579f
C318 VDD a_10976_296# 6.18e-19
C319 a_14894_160# a_15162_730# 0.030392f
C320 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15578_1376# 0.100263f
C321 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.018644f
C322 a_17176_160# a_17444_730# 0.030392f
C323 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17860_1376# 0.100263f
C324 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 6.79e-20
C325 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_4168_1376# 0.100263f
C326 a_10598_730# a_10598_296# 0.003413f
C327 a_12880_730# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 1.47e-19
C328 VDD stop 0.192279f
C329 start_buffer_0.start_delay a_n8778_3464# 1.56e-19
C330 VDD a_8694_296# 6.18e-19
C331 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 0.871529f
C332 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_12612_160# 6.08e-20
C333 a_6412_730# a_6450_1376# 0.030083f
C334 a_n8198_3464# a_n7908_3464# 0.083149f
C335 a_10330_160# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.164402f
C336 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.747722f
C337 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.010157f
C338 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 1.17e-19
C339 a_11014_1376# a_10976_730# 0.030083f
C340 VDD vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.57087f
C341 a_3752_296# a_3484_160# 1.02e-19
C342 VDD vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 3.23801f
C343 a_12880_296# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.010872f
C344 term_5 a_13296_1376# 0.014823f
C345 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1886_1376# 0.100263f
C346 a_8016_2192# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.09966f
C347 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8694_730# 0.504416f
C348 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VDD 5.07265f
C349 a_17860_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 2.36e-21
C350 a_13296_1376# a_14894_160# 0.005973f
C351 a_17176_160# VDD 1.42789f
C352 term_4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.229061f
C353 term_7 a_15578_1376# 6.12e-20
C354 VDD vernier_delay_line_0.delay_unit_2_0.out_1 2.23953f
C355 a_15162_296# a_14894_160# 1.02e-19
C356 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.001059f
C357 vernier_delay_line_0.start_neg vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.626611f
C358 term_4 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 3.69e-19
C359 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_3484_160# 1.15e-21
C360 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.019931f
C361 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 1.24e-19
C362 a_1170_2192# a_1202_160# 2.08e-21
C363 a_12880_730# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.035356f
C364 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 0.752988f
C365 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.501329f
C366 a_5766_160# term_2 0.098219f
C367 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 3.6e-19
C368 a_15162_730# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.035356f
C369 term_5 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 6.28e-22
C370 term_6 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 3.69e-19
C371 term_5 a_11014_1376# 6.12e-20
C372 a_11014_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.197073f
C373 VDD vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.706518f
C374 a_8316_730# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.003664f
C375 VDD vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.706518f
C376 term_7 a_17444_730# 0.492009f
C377 a_14894_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.164402f
C378 a_8694_730# VDD 0.497547f
C379 a_6450_1376# term_3 6.12e-20
C380 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.441403f
C381 VDD vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.706489f
C382 a_6034_296# a_6034_730# 0.003413f
C383 a_n7908_3464# a_n7618_3464# 0.083149f
C384 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 1.24e-19
C385 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_5766_160# 3.45e-19
C386 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.006183f
C387 a_1848_296# a_1848_730# 0.003413f
C388 VDD a_n8488_3464# 1.1544f
C389 a_6412_296# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.174293f
C390 vernier_delay_line_0.start_neg vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.007279f
C391 a_10298_2192# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.192064f
C392 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_6450_1376# 0.197073f
C393 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.283838f
C394 a_8048_160# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.196688f
C395 a_13296_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 7.19e-22
C396 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.001059f
C397 VDD a_12612_160# 1.42789f
C398 term_7 VDD 0.587468f
C399 a_15162_296# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.010872f
C400 a_3452_2192# a_3484_160# 2.08e-21
C401 a_8732_1376# term_3 0.014823f
C402 a_12612_160# a_12880_296# 1.02e-19
C403 a_8732_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 3.26e-19
C404 term_6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 0.229061f
C405 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 term_2 0.201251f
C406 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.132512f
C407 a_13296_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.197073f
C408 term_4 VDD 0.587468f
C409 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 3.6e-19
C410 VDD vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 3.23801f
C411 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_1 0.10528f
C412 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1848_296# 0.012202f
C413 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_6034_730# 1.47e-19
C414 a_8316_296# term_3 0.188081f
C415 term_0 a_1470_730# 0.492009f
C416 a_15540_730# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.003607f
C417 a_12612_160# a_12880_730# 0.030392f
C418 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13296_1376# 0.100263f
C419 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 0.871529f
C420 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 3.6e-19
C421 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 4.28924f
C422 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.018644f
C423 term_7 a_17822_730# 0.013457f
C424 a_17176_160# a_17444_296# 1.02e-19
C425 a_12612_160# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.45e-19
C426 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.59e-20
C427 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 3.6e-19
C428 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 a_5766_160# 4.55e-19
C429 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 3.6e-19
C430 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_1470_730# 0.035356f
C431 a_17176_160# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.164402f
C432 a_n7618_3464# a_n7328_3464# 0.083149f
C433 a_n8198_3464# a_n6748_3464# 1.76e-19
C434 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq term_2 0.229061f
C435 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 1.17e-19
C436 VDD a_n7908_3464# 1.15434f
C437 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 1.99e-19
C438 a_4168_1376# term_2 6.12e-20
C439 a_11014_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 3.26e-19
C440 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.138536f
C441 a_6412_296# VDD 6.18e-19
C442 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.953579f
C443 a_5766_160# a_6450_1376# 0.005826f
C444 term_4 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.201251f
C445 a_10330_160# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq 0.01482f
C446 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.006183f
C447 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 2.59e-20
C448 a_10330_160# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 4.55e-19
C449 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_4168_1376# 0.162625f
C450 a_8694_296# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.012202f
C451 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.132512f
C452 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 a_1886_1376# 7.19e-22
C453 a_8048_160# a_6450_1376# 0.005973f
C454 a_4130_296# a_4130_730# 0.003413f
C455 vernier_delay_line_0.start_pos vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.754929f
C456 a_17860_1376# VDD 1.40742f
C457 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.237663f
C458 term_4 a_10598_730# 0.492009f
C459 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 term_0 1.13e-20
C460 a_14862_2192# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.09966f
C461 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 7.03e-19
C462 a_15162_730# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 1.47e-19
C463 diff_gen_0.delay_unit_2_1.in_1 diff_gen_0.delay_unit_2_3.in_1 0.001356f
C464 a_8016_2192# vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.007929f
C465 a_1470_296# term_0 0.188081f
C466 a_10298_2192# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.09966f
C467 term_7 a_17444_296# 0.188081f
C468 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17822_296# 0.174293f
C469 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_10330_160# 6.08e-20
C470 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 9.61e-20
C471 term_5 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 3.69e-19
C472 a_6412_730# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.033952f
C473 term_5 a_13258_730# 0.013457f
C474 term_7 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.10528f
C475 a_8048_160# a_8732_1376# 0.005826f
C476 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_6450_1376# 0.162625f
C477 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 0.003768f
C478 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.441403f
C479 term_0 a_1848_730# 0.013457f
C480 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_11014_1376# 0.100263f
C481 a_n7618_3464# a_n6748_3464# 4.98e-19
C482 a_n7328_3464# a_n7038_3464# 0.083149f
C483 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.501329f
C484 start_buffer_0.start_delay VDD 4.0504f
C485 VDD term_2 0.587468f
C486 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.283838f
C487 diff_gen_0.delay_unit_2_1.in_1 a_n7618_3464# 2.18e-19
C488 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.237663f
C489 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.501329f
C490 VDD a_n7328_3464# 1.15434f
C491 a_10976_730# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.033952f
C492 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_1470_296# 0.010872f
C493 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.752988f
C494 a_11014_1376# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 5.04e-20
C495 VDD vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 2.57087f
C496 VDD a_15162_730# 0.497771f
C497 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq term_1 0.229061f
C498 VDD a_3752_730# 0.497771f
C499 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 1.24e-19
C500 a_15578_1376# a_15540_730# 0.030083f
C501 start_buffer_0.start_buff a_n8488_3464# 1.66e-19
C502 a_17860_1376# a_17822_730# 0.030083f
C503 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_1848_730# 0.003607f
C504 a_15578_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.197073f
C505 a_8048_160# a_8316_296# 1.02e-19
C506 a_8732_1376# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 2.36e-21
C507 VDD vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 2.57087f
C508 VDD a_1470_730# 0.497771f
C509 vernier_delay_line_0.start_pos vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 7.03e-19
C510 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 a_15578_1376# 7.19e-22
C511 a_8694_730# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.033952f
C512 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq a_6450_1376# 0.100263f
C513 a_10330_160# VDD 1.42789f
C514 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.231672f
C515 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 7.03e-19
C516 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 term_0 0.10528f
C517 a_12580_2192# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 0.192064f
C518 VDD a_13296_1376# 1.40782f
C519 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_3752_730# 1.47e-19
C520 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 term_3 6.28e-22
C521 a_15162_296# VDD 6.18e-19
C522 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 1.17e-19
C523 a_15540_296# a_15578_1376# 1.02e-19
C524 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.501329f
C525 term_5 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 1.53e-22
C526 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 3.6e-19
C527 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 term_3 1.53e-22
C528 term_6 a_15162_730# 0.492009f
C529 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.138536f
C530 term_4 a_10598_296# 0.188081f
C531 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.28924f
C532 a_1886_1376# a_1848_730# 0.030083f
C533 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.006183f
C534 a_17444_730# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.035356f
C535 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.019931f
C536 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 4.73e-19
C537 a_n7038_3464# a_n6748_3464# 0.087529f
C538 diff_gen_0.delay_unit_2_1.in_1 a_n7038_3464# 8.59e-20
C539 VDD a_n6748_3464# 1.86061f
C540 term_4 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.53e-22
C541 a_1202_160# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq 0.01482f
C542 diff_gen_0.delay_unit_2_1.in_1 VDD 4.44047f
C543 a_10330_160# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.196688f
C544 a_12612_160# vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 3.84e-19
C545 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.441403f
C546 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 a_5734_2192# 0.192064f
C547 VDD a_15540_730# 0.497547f
C548 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.283838f
C549 VDD vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 2.43248f
C550 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VDD 3.23801f
C551 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 0.441403f
C552 VDD a_11014_1376# 1.40782f
C553 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8732_1376# 0.100263f
C554 a_13296_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 2.36e-21
C555 a_12580_2192# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 1.06381f
C556 term_6 a_13296_1376# 6.12e-20
C557 a_13258_730# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.033952f
C558 a_8694_730# a_8694_296# 0.003413f
C559 term_6 a_15162_296# 0.188081f
C560 a_8016_2192# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 1.06381f
C561 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.001059f
C562 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VDD 2.55554f
C563 a_17860_1376# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.197073f
C564 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 2.59e-20
C565 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 1.24e-19
C566 vernier_delay_line_0.start_neg vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.019727f
C567 a_6034_730# term_2 0.492009f
C568 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 1.24e-19
C569 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 a_1886_1376# 0.197073f
C570 VDD vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 5.20486f
C571 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_13258_730# 0.504416f
C572 VDD a_6450_1376# 1.40782f
C573 VDD a_1470_296# 6.18e-19
C574 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.953579f
C575 a_17176_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq 6.08e-20
C576 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 a_3484_160# 3.45e-19
C577 a_10330_160# a_10598_730# 0.030392f
C578 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq a_8316_296# 0.005542f
C579 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 term_3 1.13e-20
C580 a_6412_730# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.003607f
C581 VDD a_1848_730# 0.497547f
C582 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 0.283838f
C583 a_15540_296# VDD 6.18e-19
C584 a_13296_1376# a_13258_296# 1.02e-19
C585 VDD vernier_delay_line_0.delay_unit_2_0.out_2 1.93357f
C586 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 7.03e-19
C587 term_6 a_15540_730# 0.013457f
C588 vernier_delay_line_0.start_pos vernier_delay_line_0.start_neg 0.688629f
C589 term_4 a_10976_296# 0.005542f
C590 a_12612_160# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.196688f
C591 term_6 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.10528f
C592 a_11014_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.162625f
C593 a_3752_296# VDD 6.18e-19
C594 a_8732_1376# VDD 1.40782f
C595 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.752988f
C596 a_4168_1376# a_4130_730# 0.030083f
C597 a_8316_730# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.035356f
C598 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.003768f
C599 a_17822_730# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.003607f
C600 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 9.61e-20
C601 a_14894_160# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.196688f
C602 VDD start 0.192218f
C603 term_7 a_17176_160# 0.098219f
C604 a_4168_1376# a_3484_160# 0.005826f
C605 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_5766_160# 0.164402f
C606 term_5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.10528f
C607 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.99e-19
C608 a_10298_2192# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.007929f
C609 a_8048_160# term_3 0.098219f
C610 start_buffer_0.start_buff start_buffer_0.start_delay 1.12095f
C611 a_6412_730# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.504416f
C612 a_1886_1376# a_3484_160# 0.005973f
C613 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.019931f
C614 VDD vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 2.43941f
C615 VDD a_8316_296# 6.18e-19
C616 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq a_10976_730# 0.504416f
C617 a_14894_160# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 1.15e-21
C618 a_n11872_5654# VDD 1.85997f
C619 term_6 a_15540_296# 0.005542f
C620 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 0.283838f
C621 term_5 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq 0.229061f
C622 a_1170_2192# vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 0.192064f
C623 a_12580_2192# a_12612_160# 2.08e-21
C624 a_1848_296# term_0 0.005542f
C625 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 2.59e-20
C626 a_8048_160# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 1.15e-21
C627 diff_gen_0.delay_unit_2_6.in_1 vernier_delay_line_0.start_neg 0.286409f
C628 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq a_14894_160# 6.08e-20
C629 a_8732_1376# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 7.19e-22
C630 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 term_2 6.28e-22
C631 a_3752_730# term_1 0.492009f
C632 VDD vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 5.07265f
C633 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.003768f
C634 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_3484_160# 4.55e-19
C635 a_17822_296# VDD 6.18e-19
C636 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.28924f
C637 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 term_2 1.53e-22
C638 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 term_1 0.201251f
C639 a_10330_160# a_10598_296# 1.02e-19
C640 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 a_3452_2192# 0.007929f
C641 VDD a_4130_730# 0.497547f
C642 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 4.28924f
C643 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 1.99e-19
C644 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 a_3752_730# 0.003664f
C645 a_17444_296# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 0.010872f
C646 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 0.871529f
C647 a_14862_2192# a_14894_160# 2.08e-21
C648 VDD a_3484_160# 1.42789f
C649 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 0.231672f
C650 a_10330_160# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 1.15e-21
C651 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 4.28924f
C652 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 4.28924f
C653 a_6034_296# term_2 0.188081f
C654 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.441403f
C655 a_1170_2192# vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 0.09966f
C656 a_6412_730# VDD 0.497547f
C657 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 6.79e-20
C658 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 0.501329f
C659 a_17822_730# a_17822_296# 0.003413f
C660 start_buffer_0.start_buff diff_gen_0.delay_unit_2_1.in_1 0.751615f
C661 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 a_8048_160# 3.84e-19
C662 VDD vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 3.23801f
C663 a_1848_296# a_1886_1376# 1.02e-19
C664 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_3484_160# 3.84e-19
C665 VDD a_13258_730# 0.497547f
C666 start_buffer_0.start_delay stop 6.15e-19
C667 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.231672f
C668 a_14894_160# a_15578_1376# 0.005826f
C669 a_17176_160# a_17860_1376# 0.005826f
C670 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 a_3452_2192# 0.192064f
C671 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq term_3 0.229061f
C672 a_1202_160# a_1470_730# 0.030392f
C673 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 a_4168_1376# 3.26e-19
C674 VDD a_10976_730# 0.497547f
C675 a_4130_296# a_4168_1376# 1.02e-19
C676 vernier_delay_line_0.start_pos vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 0.283838f
C677 VDD vernier_delay_line_0.start_neg 3.22778f
C678 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 0.010157f
C679 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 term_2 1.13e-20
C680 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 0.231672f
C681 a_10598_730# vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 1.47e-19
C682 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 term_0 3.69e-19
C683 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.018644f
C684 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 a_5766_160# 0.196688f
C685 a_14862_2192# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 1.06381f
C686 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 4.73e-19
C687 a_10298_2192# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 1.06381f
C688 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 9.61e-20
C689 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 a_17144_2192# 0.09966f
C690 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 1.17e-19
C691 a_14894_160# vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 3.84e-19
C692 a_8316_730# a_8316_296# 0.003413f
C693 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 a_6450_1376# 3.26e-19
C694 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 0.010157f
C695 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 0.237663f
C696 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 7.03e-19
C697 VDD a_1848_296# 6.18e-19
C698 VDD term_3 0.587468f
C699 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.283838f
C700 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 0.018644f
C701 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 7.03e-19
C702 a_10976_730# vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 0.003607f
C703 start_buffer_0.start_buff start 5.26e-19
C704 a_8048_160# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 3.45e-19
C705 a_13296_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 0.162625f
C706 VDD vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 2.43248f
C707 term_5 VDD 0.587468f
C708 a_3752_296# term_1 0.188081f
C709 term_5 a_12880_296# 0.188081f
C710 a_15578_1376# vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 0.162625f
C711 a_17822_296# vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 0.012202f
C712 VDD a_14894_160# 1.42789f
C713 a_5766_160# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 0.01482f
C714 diff_gen_0.delay_unit_2_3.in_1 diff_gen_0.delay_unit_2_4.in_1 0.756572f
C715 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq a_15162_730# 0.013457f
C716 a_13258_730# a_13258_296# 0.003413f
C717 VDD vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 2.43248f
C718 a_8732_1376# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 0.197073f
C719 term_7 a_17860_1376# 0.014823f
C720 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq a_17444_730# 0.013457f
C721 vernier_delay_line_0.start_pos vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 4.73e-19
C722 a_n11872_5654# start_buffer_0.start_buff 0.684455f
C723 diff_gen_0.delay_unit_2_1.in_1 stop 7.3e-20
C724 a_4130_296# VDD 6.18e-19
C725 a_4168_1376# a_5766_160# 0.005973f
C726 a_11014_1376# a_10976_296# 1.02e-19
C727 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 0.018644f
C728 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq a_3752_730# 0.013457f
C729 a_8694_730# vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 0.003607f
C730 diff_gen_0.delay_unit_2_4.in_1 diff_gen_0.delay_unit_2_6.in_1 0.001356f
C731 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 a_1202_160# 3.84e-19
C732 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq 0.001059f
C733 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq 0.132512f
C734 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 term_0 0.201251f
C735 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 term_1 1.53e-22
C736 a_1470_296# a_1202_160# 1.02e-19
C737 VDD a_n8778_3464# 1.15414f
C738 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 a_1886_1376# 5.04e-20
C739 diff_gen_0.delay_unit_2_6.in_1 vernier_delay_line_0.start_pos 0.728719f
C740 term_5 a_12880_730# 0.492009f
C741 a_8048_160# vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq 6.08e-20
C742 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq a_1470_730# 0.013457f
C743 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 0.747722f
C744 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 0.441403f
C745 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 7.03e-19
C746 a_11014_1376# vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 7.19e-22
C747 term_7 VSS 0.712334f
C748 term_6 VSS 0.712333f
C749 term_5 VSS 0.712333f
C750 term_4 VSS 0.712333f
C751 term_3 VSS 0.712333f
C752 term_2 VSS 0.712333f
C753 term_1 VSS 0.712333f
C754 term_0 VSS 0.712422f
C755 stop VSS 0.268426f
C756 start VSS 0.268973f
C757 VDD VSS 0.212509p
C758 a_17822_296# VSS 0.192129f
C759 a_17444_296# VSS 0.190624f
C760 a_15540_296# VSS 0.192129f
C761 a_17822_730# VSS 0.023462f
C762 a_15162_296# VSS 0.190624f
C763 a_17444_730# VSS 0.024712f
C764 a_17860_1376# VSS 0.830566f
C765 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nq VSS 0.583498f
C766 a_17176_160# VSS 0.829382f
C767 a_13258_296# VSS 0.192129f
C768 a_15540_730# VSS 0.023462f
C769 a_12880_296# VSS 0.190624f
C770 a_15162_730# VSS 0.024712f
C771 a_15578_1376# VSS 0.823407f
C772 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.nq VSS 0.583296f
C773 a_14894_160# VSS 0.829382f
C774 a_10976_296# VSS 0.192129f
C775 a_13258_730# VSS 0.023462f
C776 a_10598_296# VSS 0.190624f
C777 a_12880_730# VSS 0.024712f
C778 a_13296_1376# VSS 0.823407f
C779 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.nq VSS 0.583296f
C780 a_12612_160# VSS 0.829382f
C781 a_8694_296# VSS 0.192129f
C782 a_10976_730# VSS 0.023462f
C783 a_8316_296# VSS 0.190624f
C784 a_10598_730# VSS 0.024712f
C785 a_11014_1376# VSS 0.823407f
C786 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.nq VSS 0.583296f
C787 a_10330_160# VSS 0.829382f
C788 a_6412_296# VSS 0.192129f
C789 a_8694_730# VSS 0.023462f
C790 a_6034_296# VSS 0.190624f
C791 a_8316_730# VSS 0.024712f
C792 a_8732_1376# VSS 0.823407f
C793 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.nq VSS 0.583296f
C794 a_8048_160# VSS 0.829382f
C795 a_4130_296# VSS 0.192129f
C796 a_6412_730# VSS 0.023462f
C797 a_3752_296# VSS 0.190624f
C798 a_6034_730# VSS 0.024712f
C799 a_6450_1376# VSS 0.823407f
C800 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.nq VSS 0.583296f
C801 a_5766_160# VSS 0.829382f
C802 a_1848_296# VSS 0.192269f
C803 a_4130_730# VSS 0.023462f
C804 a_1470_296# VSS 0.190873f
C805 a_3752_730# VSS 0.024712f
C806 a_4168_1376# VSS 0.823407f
C807 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.nq VSS 0.583296f
C808 a_3484_160# VSS 0.829382f
C809 a_1848_730# VSS 0.023462f
C810 a_1470_730# VSS 0.024712f
C811 a_1886_1376# VSS 0.82359f
C812 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.nq VSS 0.583876f
C813 a_1202_160# VSS 0.838649f
C814 a_17144_2192# VSS 0.354057f
C815 a_14862_2192# VSS 0.354057f
C816 a_12580_2192# VSS 0.354057f
C817 a_10298_2192# VSS 0.354057f
C818 a_8016_2192# VSS 0.354057f
C819 a_5734_2192# VSS 0.354057f
C820 a_3452_2192# VSS 0.354057f
C821 a_1170_2192# VSS 0.354057f
C822 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1 VSS 6.49614f
C823 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2 VSS 6.442006f
C824 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C825 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C826 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C827 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C828 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C829 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C830 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C831 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C832 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C833 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C834 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1 VSS 6.023691f
C835 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2 VSS 6.442516f
C836 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1 VSS 6.025101f
C837 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2 VSS 7.090996f
C838 a_n6748_3464# VSS 1.4918f
C839 a_n7038_3464# VSS 0.622536f
C840 a_n7328_3464# VSS 0.622289f
C841 a_n7618_3464# VSS 0.622523f
C842 a_n7908_3464# VSS 0.622248f
C843 a_n8198_3464# VSS 0.622523f
C844 a_n8488_3464# VSS 0.622523f
C845 a_n8778_3464# VSS 0.630914f
C846 vernier_delay_line_0.delay_unit_2_0.out_2 VSS 1.24637f
C847 vernier_delay_line_0.delay_unit_2_0.out_1 VSS 0.974288f
C848 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2 VSS 6.020628f
C849 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1 VSS 5.680524f
C850 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2 VSS 6.071241f
C851 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1 VSS 5.680524f
C852 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2 VSS 6.071241f
C853 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1 VSS 5.488731f
C854 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2 VSS 6.071241f
C855 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1 VSS 5.488731f
C856 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2 VSS 6.071241f
C857 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1 VSS 5.680524f
C858 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2 VSS 6.020628f
C859 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1 VSS 5.680524f
C860 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2 VSS 6.020728f
C861 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1 VSS 5.655783f
C862 vernier_delay_line_0.start_neg VSS 3.59562f
C863 vernier_delay_line_0.start_pos VSS 2.779078f
C864 diff_gen_0.delay_unit_2_6.in_1 VSS 2.070971f
C865 diff_gen_0.delay_unit_2_4.in_1 VSS 2.006581f
C866 diff_gen_0.delay_unit_2_3.in_1 VSS 2.006331f
C867 diff_gen_0.delay_unit_2_1.in_1 VSS 2.012701f
C868 start_buffer_0.start_delay VSS 3.817548f
C869 start_buffer_0.start_buff VSS 5.282834f
C870 a_n11872_5654# VSS 1.50746f
C871 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.936187f
C872 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.087567f
C873 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.039891f
C874 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.097546f
C875 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C876 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C877 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C878 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.115133f
C879 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.095888f
C880 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.041221f
C881 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C882 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.108538f
C883 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.081767f
C884 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.090596f
C885 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C886 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C887 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.398296f
C888 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.36504f
C889 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out2.n7 VSS 0.753756f
C890 a_17320_2192.t1 VSS 0.059028f
C891 a_17320_2192.t5 VSS 0.059028f
C892 a_17320_2192.t4 VSS 0.059028f
C893 a_17320_2192.n0 VSS 0.139449f
C894 a_17320_2192.t2 VSS 0.059028f
C895 a_17320_2192.t0 VSS 0.059028f
C896 a_17320_2192.n1 VSS 0.136068f
C897 a_17320_2192.n2 VSS 1.11221f
C898 a_17320_2192.n3 VSS 0.258102f
C899 a_17320_2192.t3 VSS 0.059028f
C900 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C901 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.096169f
C902 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.041341f
C903 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.116331f
C904 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C905 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C906 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.114315f
C907 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.202807f
C908 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.087824f
C909 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.040008f
C910 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.097717f
C911 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.200111f
C912 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.382243f
C913 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.107599f
C914 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C915 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.082007f
C916 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.090862f
C917 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.108213f
C918 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.out1.n7 VSS 1.24645f
C919 a_1346_2192.t2 VSS 0.059028f
C920 a_1346_2192.t0 VSS 0.059028f
C921 a_1346_2192.t1 VSS 0.059028f
C922 a_1346_2192.n0 VSS 0.139449f
C923 a_1346_2192.t3 VSS 0.059028f
C924 a_1346_2192.t5 VSS 0.059028f
C925 a_1346_2192.n1 VSS 0.258102f
C926 a_1346_2192.n2 VSS 1.11221f
C927 a_1346_2192.n3 VSS 0.136068f
C928 a_1346_2192.t4 VSS 0.059028f
C929 a_3628_2192.t1 VSS 0.059028f
C930 a_3628_2192.t5 VSS 0.059028f
C931 a_3628_2192.t4 VSS 0.059028f
C932 a_3628_2192.n0 VSS 0.139449f
C933 a_3628_2192.t2 VSS 0.059028f
C934 a_3628_2192.t0 VSS 0.059028f
C935 a_3628_2192.n1 VSS 0.136068f
C936 a_3628_2192.n2 VSS 1.11221f
C937 a_3628_2192.n3 VSS 0.258102f
C938 a_3628_2192.t3 VSS 0.059028f
C939 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.936187f
C940 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.087567f
C941 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.039891f
C942 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.097546f
C943 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C944 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C945 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C946 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.115133f
C947 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.095888f
C948 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.041221f
C949 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C950 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.108538f
C951 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.081767f
C952 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.090596f
C953 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C954 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C955 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.398296f
C956 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.36504f
C957 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out2.n7 VSS 0.753756f
C958 vernier_delay_line_0.delay_unit_2_0.out_1.t2 VSS 0.020532f
C959 vernier_delay_line_0.delay_unit_2_0.out_1.t1 VSS 0.020532f
C960 vernier_delay_line_0.delay_unit_2_0.out_1.n0 VSS 0.048092f
C961 vernier_delay_line_0.delay_unit_2_0.out_1.t3 VSS 0.061597f
C962 vernier_delay_line_0.delay_unit_2_0.out_1.t5 VSS 0.061597f
C963 vernier_delay_line_0.delay_unit_2_0.out_1.n1 VSS 0.125485f
C964 vernier_delay_line_0.delay_unit_2_0.out_1.n2 VSS 0.522094f
C965 vernier_delay_line_0.delay_unit_2_0.out_1.t0 VSS 0.075157f
C966 vernier_delay_line_0.delay_unit_2_0.out_1.t4 VSS 0.227425f
C967 vernier_delay_line_0.delay_unit_2_0.out_1.n3 VSS 0.55466f
C968 vernier_delay_line_0.delay_unit_2_0.out_1.n4 VSS 0.283681f
C969 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C970 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.096169f
C971 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.041341f
C972 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.116331f
C973 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C974 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C975 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.114315f
C976 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.202807f
C977 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.087824f
C978 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.040008f
C979 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.097717f
C980 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.200111f
C981 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.382243f
C982 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.107599f
C983 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C984 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.082007f
C985 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.090862f
C986 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.108213f
C987 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.out1.n7 VSS 1.24645f
C988 diff_gen_0.delay_unit_2_4.in_2.t10 VSS 0.066664f
C989 diff_gen_0.delay_unit_2_4.in_2.t13 VSS 0.021266f
C990 diff_gen_0.delay_unit_2_4.in_2.n0 VSS 0.046756f
C991 diff_gen_0.delay_unit_2_4.in_2.t15 VSS 0.066664f
C992 diff_gen_0.delay_unit_2_4.in_2.t9 VSS 0.021266f
C993 diff_gen_0.delay_unit_2_4.in_2.n1 VSS 0.046454f
C994 diff_gen_0.delay_unit_2_4.in_2.n2 VSS 0.014982f
C995 diff_gen_0.delay_unit_2_4.in_2.t12 VSS 0.066664f
C996 diff_gen_0.delay_unit_2_4.in_2.t14 VSS 0.021266f
C997 diff_gen_0.delay_unit_2_4.in_2.n3 VSS 0.046756f
C998 diff_gen_0.delay_unit_2_4.in_2.t8 VSS 0.066664f
C999 diff_gen_0.delay_unit_2_4.in_2.t11 VSS 0.021266f
C1000 diff_gen_0.delay_unit_2_4.in_2.n4 VSS 0.046454f
C1001 diff_gen_0.delay_unit_2_4.in_2.n5 VSS 0.014821f
C1002 diff_gen_0.delay_unit_2_4.in_2.n6 VSS 0.22891f
C1003 diff_gen_0.delay_unit_2_4.in_2.t7 VSS 0.165681f
C1004 diff_gen_0.delay_unit_2_4.in_2.t6 VSS 0.051203f
C1005 diff_gen_0.delay_unit_2_4.in_2.n7 VSS 0.452839f
C1006 diff_gen_0.delay_unit_2_4.in_2.n8 VSS 0.285821f
C1007 diff_gen_0.delay_unit_2_4.in_2.t3 VSS 0.043739f
C1008 diff_gen_0.delay_unit_2_4.in_2.t4 VSS 0.043739f
C1009 diff_gen_0.delay_unit_2_4.in_2.n9 VSS 0.093535f
C1010 diff_gen_0.delay_unit_2_4.in_2.t2 VSS 0.01458f
C1011 diff_gen_0.delay_unit_2_4.in_2.t0 VSS 0.01458f
C1012 diff_gen_0.delay_unit_2_4.in_2.n10 VSS 0.031652f
C1013 diff_gen_0.delay_unit_2_4.in_2.n11 VSS 0.376142f
C1014 diff_gen_0.delay_unit_2_4.in_2.t5 VSS 0.165681f
C1015 diff_gen_0.delay_unit_2_4.in_2.t1 VSS 0.051203f
C1016 diff_gen_0.delay_unit_2_4.in_2.n12 VSS 0.398173f
C1017 diff_gen_0.delay_unit_2_4.in_2.n13 VSS 0.085944f
C1018 diff_gen_0.delay_unit_2_3.out_2 VSS 0.028637f
C1019 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.096169f
C1020 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.041341f
C1021 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C1022 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C1023 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1024 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C1025 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.202807f
C1026 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.087824f
C1027 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.040008f
C1028 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C1029 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C1030 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C1031 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C1032 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C1033 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.107599f
C1034 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C1035 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.082007f
C1036 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.090862f
C1037 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C1038 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C1039 a_12756_2192.t1 VSS 0.059028f
C1040 a_12756_2192.t4 VSS 0.059028f
C1041 a_12756_2192.t5 VSS 0.059028f
C1042 a_12756_2192.n0 VSS 0.139449f
C1043 a_12756_2192.t0 VSS 0.059028f
C1044 a_12756_2192.t2 VSS 0.059028f
C1045 a_12756_2192.n1 VSS 0.136068f
C1046 a_12756_2192.n2 VSS 1.11221f
C1047 a_12756_2192.n3 VSS 0.258102f
C1048 a_12756_2192.t3 VSS 0.059028f
C1049 a_8192_2192.t2 VSS 0.059028f
C1050 a_8192_2192.t1 VSS 0.059028f
C1051 a_8192_2192.t0 VSS 0.059028f
C1052 a_8192_2192.n0 VSS 0.139449f
C1053 a_8192_2192.t5 VSS 0.059028f
C1054 a_8192_2192.t3 VSS 0.059028f
C1055 a_8192_2192.n1 VSS 0.258102f
C1056 a_8192_2192.n2 VSS 1.11221f
C1057 a_8192_2192.n3 VSS 0.136068f
C1058 a_8192_2192.t4 VSS 0.059028f
C1059 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.096169f
C1060 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.041341f
C1061 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C1062 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C1063 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1064 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C1065 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.202807f
C1066 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.087824f
C1067 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.040008f
C1068 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C1069 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.200111f
C1070 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C1071 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C1072 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C1073 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.107599f
C1074 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C1075 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.082007f
C1076 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.090862f
C1077 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C1078 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C1079 a_10210_2192.t10 VSS 0.024913f
C1080 a_10210_2192.t12 VSS 0.024913f
C1081 a_10210_2192.t9 VSS 0.024913f
C1082 a_10210_2192.n0 VSS 0.057409f
C1083 a_10210_2192.t0 VSS 0.024913f
C1084 a_10210_2192.t4 VSS 0.024913f
C1085 a_10210_2192.n1 VSS 0.060114f
C1086 a_10210_2192.t6 VSS 0.024913f
C1087 a_10210_2192.t3 VSS 0.024913f
C1088 a_10210_2192.n2 VSS 0.060114f
C1089 a_10210_2192.t1 VSS 0.024913f
C1090 a_10210_2192.t5 VSS 0.024913f
C1091 a_10210_2192.n3 VSS 0.060114f
C1092 a_10210_2192.t7 VSS 0.097139f
C1093 a_10210_2192.n4 VSS 0.369186f
C1094 a_10210_2192.n5 VSS 0.182473f
C1095 a_10210_2192.n6 VSS 0.22019f
C1096 a_10210_2192.t8 VSS 0.024913f
C1097 a_10210_2192.t2 VSS 0.024913f
C1098 a_10210_2192.n7 VSS 0.052659f
C1099 a_10210_2192.n8 VSS 0.140942f
C1100 a_10210_2192.n9 VSS 0.340434f
C1101 a_10210_2192.n10 VSS 0.060272f
C1102 a_10210_2192.t11 VSS 0.024913f
C1103 a_10474_2192.t5 VSS 0.059028f
C1104 a_10474_2192.t3 VSS 0.059028f
C1105 a_10474_2192.t0 VSS 0.059028f
C1106 a_10474_2192.n0 VSS 0.136068f
C1107 a_10474_2192.t2 VSS 0.059028f
C1108 a_10474_2192.t1 VSS 0.059028f
C1109 a_10474_2192.n1 VSS 0.258102f
C1110 a_10474_2192.n2 VSS 1.11221f
C1111 a_10474_2192.n3 VSS 0.139449f
C1112 a_10474_2192.t4 VSS 0.059028f
C1113 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t10 VSS 0.039259f
C1114 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t12 VSS 0.012524f
C1115 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n0 VSS 0.027534f
C1116 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t16 VSS 0.039259f
C1117 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t19 VSS 0.012524f
C1118 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1119 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1120 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t8 VSS 0.039259f
C1121 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t11 VSS 0.012524f
C1122 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n3 VSS 0.027534f
C1123 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t14 VSS 0.039259f
C1124 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t17 VSS 0.012524f
C1125 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1126 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1127 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1128 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t1 VSS 0.09757f
C1129 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t0 VSS 0.030153f
C1130 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1131 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t9 VSS 0.046129f
C1132 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t15 VSS 0.046129f
C1133 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1134 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t13 VSS 0.046129f
C1135 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t18 VSS 0.046129f
C1136 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1137 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1138 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t7 VSS 0.025758f
C1139 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t6 VSS 0.025758f
C1140 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1141 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t3 VSS 0.008586f
C1142 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t2 VSS 0.008586f
C1143 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1144 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1145 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t5 VSS 0.09757f
C1146 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.t4 VSS 0.030153f
C1147 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1148 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n15 VSS 0.050613f
C1149 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_2.n16 VSS 0.122976f
C1150 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.096169f
C1151 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.041341f
C1152 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n0 VSS 0.116331f
C1153 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C1154 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1155 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.114315f
C1156 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.202807f
C1157 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.087824f
C1158 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.040008f
C1159 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.097717f
C1160 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C1161 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.661409f
C1162 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.399989f
C1163 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.382243f
C1164 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.107599f
C1165 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.139678f
C1166 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.082007f
C1167 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.090862f
C1168 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.108213f
C1169 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out1.n8 VSS 1.24645f
C1170 a_17056_2192.t10 VSS 0.024913f
C1171 a_17056_2192.t9 VSS 0.024913f
C1172 a_17056_2192.t12 VSS 0.024913f
C1173 a_17056_2192.n0 VSS 0.060272f
C1174 a_17056_2192.t4 VSS 0.024913f
C1175 a_17056_2192.t2 VSS 0.024913f
C1176 a_17056_2192.n1 VSS 0.060114f
C1177 a_17056_2192.t0 VSS 0.024913f
C1178 a_17056_2192.t6 VSS 0.024913f
C1179 a_17056_2192.n2 VSS 0.060114f
C1180 a_17056_2192.t7 VSS 0.024913f
C1181 a_17056_2192.t3 VSS 0.024913f
C1182 a_17056_2192.n3 VSS 0.060114f
C1183 a_17056_2192.t1 VSS 0.097139f
C1184 a_17056_2192.n4 VSS 0.369186f
C1185 a_17056_2192.n5 VSS 0.182473f
C1186 a_17056_2192.n6 VSS 0.22019f
C1187 a_17056_2192.t8 VSS 0.024913f
C1188 a_17056_2192.t5 VSS 0.024913f
C1189 a_17056_2192.n7 VSS 0.052659f
C1190 a_17056_2192.n8 VSS 0.140942f
C1191 a_17056_2192.n9 VSS 0.340434f
C1192 a_17056_2192.n10 VSS 0.057409f
C1193 a_17056_2192.t11 VSS 0.024913f
C1194 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t18 VSS 0.061029f
C1195 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t8 VSS 0.019469f
C1196 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n0 VSS 0.042527f
C1197 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t11 VSS 0.061029f
C1198 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t14 VSS 0.019469f
C1199 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n1 VSS 0.042803f
C1200 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n2 VSS 0.013718f
C1201 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t17 VSS 0.061029f
C1202 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t19 VSS 0.019469f
C1203 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n3 VSS 0.042803f
C1204 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t9 VSS 0.061029f
C1205 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t13 VSS 0.019469f
C1206 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n4 VSS 0.042527f
C1207 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n5 VSS 0.013568f
C1208 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n6 VSS 0.358094f
C1209 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t6 VSS 0.048842f
C1210 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t7 VSS 0.14784f
C1211 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n7 VSS 0.375222f
C1212 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n8 VSS 0.195554f
C1213 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t2 VSS 0.013347f
C1214 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t1 VSS 0.013347f
C1215 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n9 VSS 0.031263f
C1216 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t5 VSS 0.040042f
C1217 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t4 VSS 0.040042f
C1218 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n10 VSS 0.081573f
C1219 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n11 VSS 0.339393f
C1220 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t10 VSS 0.062678f
C1221 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t15 VSS 0.062678f
C1222 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n12 VSS 0.070759f
C1223 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t16 VSS 0.062678f
C1224 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t12 VSS 0.062678f
C1225 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n13 VSS 0.070376f
C1226 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n14 VSS 0.642547f
C1227 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t0 VSS 0.046875f
C1228 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n15 VSS 0.161895f
C1229 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.t3 VSS 0.14784f
C1230 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n16 VSS 0.245357f
C1231 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_1.n17 VSS 0.18441f
C1232 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1233 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1234 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.087567f
C1235 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.039891f
C1236 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1237 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1238 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C1239 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C1240 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.115133f
C1241 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.095888f
C1242 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.041221f
C1243 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.116123f
C1244 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.108538f
C1245 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.081767f
C1246 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.090596f
C1247 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.106694f
C1248 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C1249 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1250 diff_gen_0.delay_unit_2_3.in_1.t11 VSS 0.086195f
C1251 diff_gen_0.delay_unit_2_3.in_1.t13 VSS 0.027496f
C1252 diff_gen_0.delay_unit_2_3.in_1.n0 VSS 0.060063f
C1253 diff_gen_0.delay_unit_2_3.in_1.t15 VSS 0.086195f
C1254 diff_gen_0.delay_unit_2_3.in_1.t9 VSS 0.027496f
C1255 diff_gen_0.delay_unit_2_3.in_1.n1 VSS 0.060453f
C1256 diff_gen_0.delay_unit_2_3.in_1.n2 VSS 0.019374f
C1257 diff_gen_0.delay_unit_2_3.in_1.t12 VSS 0.086195f
C1258 diff_gen_0.delay_unit_2_3.in_1.t14 VSS 0.027496f
C1259 diff_gen_0.delay_unit_2_3.in_1.n3 VSS 0.060453f
C1260 diff_gen_0.delay_unit_2_3.in_1.t8 VSS 0.086195f
C1261 diff_gen_0.delay_unit_2_3.in_1.t10 VSS 0.027496f
C1262 diff_gen_0.delay_unit_2_3.in_1.n4 VSS 0.060063f
C1263 diff_gen_0.delay_unit_2_3.in_1.n5 VSS 0.019163f
C1264 diff_gen_0.delay_unit_2_3.in_1.n6 VSS 0.505752f
C1265 diff_gen_0.delay_unit_2_3.in_1.t6 VSS 0.068982f
C1266 diff_gen_0.delay_unit_2_3.in_1.t7 VSS 0.2088f
C1267 diff_gen_0.delay_unit_2_3.in_1.n7 VSS 0.529943f
C1268 diff_gen_0.delay_unit_2_3.in_1.n8 VSS 0.27619f
C1269 diff_gen_0.delay_unit_2_3.in_1.t2 VSS 0.018851f
C1270 diff_gen_0.delay_unit_2_3.in_1.t0 VSS 0.018851f
C1271 diff_gen_0.delay_unit_2_3.in_1.n9 VSS 0.044154f
C1272 diff_gen_0.delay_unit_2_3.in_1.t5 VSS 0.056553f
C1273 diff_gen_0.delay_unit_2_3.in_1.t3 VSS 0.056553f
C1274 diff_gen_0.delay_unit_2_3.in_1.n10 VSS 0.115209f
C1275 diff_gen_0.delay_unit_2_3.in_1.n11 VSS 0.479339f
C1276 diff_gen_0.delay_unit_2_3.in_1.t1 VSS 0.069002f
C1277 diff_gen_0.delay_unit_2_3.in_1.t4 VSS 0.2088f
C1278 diff_gen_0.delay_unit_2_3.in_1.n12 VSS 0.509237f
C1279 diff_gen_0.delay_unit_2_3.in_1.n13 VSS 0.26045f
C1280 diff_gen_0.delay_unit_2_2.in_2.t10 VSS 0.066664f
C1281 diff_gen_0.delay_unit_2_2.in_2.t12 VSS 0.021266f
C1282 diff_gen_0.delay_unit_2_2.in_2.n0 VSS 0.046756f
C1283 diff_gen_0.delay_unit_2_2.in_2.t8 VSS 0.066664f
C1284 diff_gen_0.delay_unit_2_2.in_2.t11 VSS 0.021266f
C1285 diff_gen_0.delay_unit_2_2.in_2.n1 VSS 0.046454f
C1286 diff_gen_0.delay_unit_2_2.in_2.n2 VSS 0.014982f
C1287 diff_gen_0.delay_unit_2_2.in_2.t13 VSS 0.066664f
C1288 diff_gen_0.delay_unit_2_2.in_2.t14 VSS 0.021266f
C1289 diff_gen_0.delay_unit_2_2.in_2.n3 VSS 0.046756f
C1290 diff_gen_0.delay_unit_2_2.in_2.t15 VSS 0.066664f
C1291 diff_gen_0.delay_unit_2_2.in_2.t9 VSS 0.021266f
C1292 diff_gen_0.delay_unit_2_2.in_2.n4 VSS 0.046454f
C1293 diff_gen_0.delay_unit_2_2.in_2.n5 VSS 0.014821f
C1294 diff_gen_0.delay_unit_2_2.in_2.n6 VSS 0.22891f
C1295 diff_gen_0.delay_unit_2_2.in_2.t1 VSS 0.165681f
C1296 diff_gen_0.delay_unit_2_2.in_2.t0 VSS 0.051203f
C1297 diff_gen_0.delay_unit_2_2.in_2.n7 VSS 0.452839f
C1298 diff_gen_0.delay_unit_2_2.in_2.n8 VSS 0.285821f
C1299 diff_gen_0.delay_unit_2_2.in_2.t5 VSS 0.043739f
C1300 diff_gen_0.delay_unit_2_2.in_2.t6 VSS 0.043739f
C1301 diff_gen_0.delay_unit_2_2.in_2.n9 VSS 0.093535f
C1302 diff_gen_0.delay_unit_2_2.in_2.t4 VSS 0.01458f
C1303 diff_gen_0.delay_unit_2_2.in_2.t2 VSS 0.01458f
C1304 diff_gen_0.delay_unit_2_2.in_2.n10 VSS 0.031652f
C1305 diff_gen_0.delay_unit_2_2.in_2.n11 VSS 0.376142f
C1306 diff_gen_0.delay_unit_2_2.in_2.t7 VSS 0.165681f
C1307 diff_gen_0.delay_unit_2_2.in_2.t3 VSS 0.051203f
C1308 diff_gen_0.delay_unit_2_2.in_2.n12 VSS 0.398173f
C1309 diff_gen_0.delay_unit_2_2.in_2.n13 VSS 0.085944f
C1310 diff_gen_0.delay_unit_2_1.out_2 VSS 0.028637f
C1311 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t17 VSS 0.059856f
C1312 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t9 VSS 0.019094f
C1313 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n0 VSS 0.041709f
C1314 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t11 VSS 0.059856f
C1315 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t14 VSS 0.019094f
C1316 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n1 VSS 0.04198f
C1317 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n2 VSS 0.013454f
C1318 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t16 VSS 0.059856f
C1319 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t8 VSS 0.019094f
C1320 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n3 VSS 0.04198f
C1321 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t10 VSS 0.059856f
C1322 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t13 VSS 0.019094f
C1323 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n4 VSS 0.041709f
C1324 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n5 VSS 0.013307f
C1325 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n6 VSS 0.351208f
C1326 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t0 VSS 0.047903f
C1327 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t1 VSS 0.144997f
C1328 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n7 VSS 0.368007f
C1329 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n8 VSS 0.191794f
C1330 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t3 VSS 0.013091f
C1331 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t2 VSS 0.013091f
C1332 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n9 VSS 0.030662f
C1333 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t7 VSS 0.039272f
C1334 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t6 VSS 0.039272f
C1335 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n10 VSS 0.080004f
C1336 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n11 VSS 0.332866f
C1337 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t19 VSS 0.061472f
C1338 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t15 VSS 0.061472f
C1339 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n12 VSS 0.069399f
C1340 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t18 VSS 0.061472f
C1341 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t12 VSS 0.061472f
C1342 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n13 VSS 0.069022f
C1343 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n14 VSS 0.63019f
C1344 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t4 VSS 0.045973f
C1345 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n15 VSS 0.158781f
C1346 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.t5 VSS 0.144997f
C1347 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n16 VSS 0.240639f
C1348 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_1.n17 VSS 0.180864f
C1349 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t17 VSS 0.039259f
C1350 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t8 VSS 0.012524f
C1351 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n0 VSS 0.027534f
C1352 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t10 VSS 0.039259f
C1353 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t13 VSS 0.012524f
C1354 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1355 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1356 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t15 VSS 0.039259f
C1357 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t18 VSS 0.012524f
C1358 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n3 VSS 0.027534f
C1359 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t11 VSS 0.039259f
C1360 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t14 VSS 0.012524f
C1361 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1362 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1363 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1364 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t0 VSS 0.09757f
C1365 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t1 VSS 0.030153f
C1366 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1367 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t16 VSS 0.046129f
C1368 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t9 VSS 0.046129f
C1369 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1370 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t19 VSS 0.046129f
C1371 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t12 VSS 0.046129f
C1372 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1373 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1374 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t7 VSS 0.025758f
C1375 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t6 VSS 0.025758f
C1376 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1377 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t4 VSS 0.008586f
C1378 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t3 VSS 0.008586f
C1379 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1380 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1381 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t5 VSS 0.09757f
C1382 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.t2 VSS 0.030153f
C1383 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1384 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n15 VSS 0.050613f
C1385 vernier_delay_line_0.saff_delay_unit_1/delay_unit_2_0.in_2.n16 VSS 0.122976f
C1386 vernier_delay_line_0.start_pos.t11 VSS 0.086445f
C1387 vernier_delay_line_0.start_pos.t13 VSS 0.027576f
C1388 vernier_delay_line_0.start_pos.n0 VSS 0.060238f
C1389 vernier_delay_line_0.start_pos.t8 VSS 0.086445f
C1390 vernier_delay_line_0.start_pos.t10 VSS 0.027576f
C1391 vernier_delay_line_0.start_pos.n1 VSS 0.060629f
C1392 vernier_delay_line_0.start_pos.n2 VSS 0.01943f
C1393 vernier_delay_line_0.start_pos.t9 VSS 0.086445f
C1394 vernier_delay_line_0.start_pos.t12 VSS 0.027576f
C1395 vernier_delay_line_0.start_pos.n3 VSS 0.060629f
C1396 vernier_delay_line_0.start_pos.t14 VSS 0.086445f
C1397 vernier_delay_line_0.start_pos.t15 VSS 0.027576f
C1398 vernier_delay_line_0.start_pos.n4 VSS 0.060238f
C1399 vernier_delay_line_0.start_pos.n5 VSS 0.019219f
C1400 vernier_delay_line_0.start_pos.n6 VSS 0.507224f
C1401 vernier_delay_line_0.start_pos.t0 VSS 0.069183f
C1402 vernier_delay_line_0.start_pos.t1 VSS 0.209408f
C1403 vernier_delay_line_0.start_pos.n7 VSS 0.531486f
C1404 vernier_delay_line_0.start_pos.n8 VSS 0.276994f
C1405 vernier_delay_line_0.start_pos.t2 VSS 0.018906f
C1406 vernier_delay_line_0.start_pos.t3 VSS 0.018906f
C1407 vernier_delay_line_0.start_pos.n9 VSS 0.044282f
C1408 vernier_delay_line_0.start_pos.t7 VSS 0.056718f
C1409 vernier_delay_line_0.start_pos.t5 VSS 0.056718f
C1410 vernier_delay_line_0.start_pos.n10 VSS 0.115544f
C1411 vernier_delay_line_0.start_pos.n11 VSS 0.480734f
C1412 vernier_delay_line_0.start_pos.t4 VSS 0.069203f
C1413 vernier_delay_line_0.start_pos.t6 VSS 0.209408f
C1414 vernier_delay_line_0.start_pos.n12 VSS 0.51072f
C1415 vernier_delay_line_0.start_pos.n13 VSS 0.261208f
C1416 a_7928_2192.t5 VSS 0.024913f
C1417 a_7928_2192.t7 VSS 0.024913f
C1418 a_7928_2192.t6 VSS 0.024913f
C1419 a_7928_2192.n0 VSS 0.060272f
C1420 a_7928_2192.t11 VSS 0.024913f
C1421 a_7928_2192.t0 VSS 0.024913f
C1422 a_7928_2192.n1 VSS 0.060114f
C1423 a_7928_2192.t2 VSS 0.024913f
C1424 a_7928_2192.t12 VSS 0.024913f
C1425 a_7928_2192.n2 VSS 0.060114f
C1426 a_7928_2192.t10 VSS 0.024913f
C1427 a_7928_2192.t1 VSS 0.024913f
C1428 a_7928_2192.n3 VSS 0.060114f
C1429 a_7928_2192.t3 VSS 0.097139f
C1430 a_7928_2192.n4 VSS 0.369186f
C1431 a_7928_2192.n5 VSS 0.182473f
C1432 a_7928_2192.n6 VSS 0.22019f
C1433 a_7928_2192.t4 VSS 0.024913f
C1434 a_7928_2192.t9 VSS 0.024913f
C1435 a_7928_2192.n7 VSS 0.052659f
C1436 a_7928_2192.n8 VSS 0.140942f
C1437 a_7928_2192.n9 VSS 0.340434f
C1438 a_7928_2192.n10 VSS 0.057409f
C1439 a_7928_2192.t8 VSS 0.024913f
C1440 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t18 VSS 0.061472f
C1441 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t10 VSS 0.061472f
C1442 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n0 VSS 0.069399f
C1443 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t13 VSS 0.061472f
C1444 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t15 VSS 0.061472f
C1445 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n1 VSS 0.069022f
C1446 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n2 VSS 0.63019f
C1447 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t14 VSS 0.059856f
C1448 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t17 VSS 0.019094f
C1449 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n3 VSS 0.041709f
C1450 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t19 VSS 0.059856f
C1451 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t9 VSS 0.019094f
C1452 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n4 VSS 0.04198f
C1453 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n5 VSS 0.013454f
C1454 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t12 VSS 0.059856f
C1455 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t16 VSS 0.019094f
C1456 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n6 VSS 0.04198f
C1457 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t8 VSS 0.059856f
C1458 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t11 VSS 0.019094f
C1459 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n7 VSS 0.041709f
C1460 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n8 VSS 0.013307f
C1461 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n9 VSS 0.351208f
C1462 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t6 VSS 0.047903f
C1463 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t7 VSS 0.144997f
C1464 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n10 VSS 0.368007f
C1465 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t1 VSS 0.013091f
C1466 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t5 VSS 0.013091f
C1467 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n11 VSS 0.030662f
C1468 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t4 VSS 0.039272f
C1469 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t3 VSS 0.039272f
C1470 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n12 VSS 0.080004f
C1471 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n13 VSS 0.332866f
C1472 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n14 VSS 0.180864f
C1473 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t0 VSS 0.144997f
C1474 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n15 VSS 0.240639f
C1475 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.t2 VSS 0.045973f
C1476 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_1.n16 VSS 0.158781f
C1477 diff_gen_0.delay_unit_2_6.in_2.t14 VSS 0.066664f
C1478 diff_gen_0.delay_unit_2_6.in_2.t8 VSS 0.021266f
C1479 diff_gen_0.delay_unit_2_6.in_2.n0 VSS 0.046756f
C1480 diff_gen_0.delay_unit_2_6.in_2.t11 VSS 0.066664f
C1481 diff_gen_0.delay_unit_2_6.in_2.t13 VSS 0.021266f
C1482 diff_gen_0.delay_unit_2_6.in_2.n1 VSS 0.046454f
C1483 diff_gen_0.delay_unit_2_6.in_2.n2 VSS 0.014982f
C1484 diff_gen_0.delay_unit_2_6.in_2.t15 VSS 0.066664f
C1485 diff_gen_0.delay_unit_2_6.in_2.t9 VSS 0.021266f
C1486 diff_gen_0.delay_unit_2_6.in_2.n3 VSS 0.046756f
C1487 diff_gen_0.delay_unit_2_6.in_2.t10 VSS 0.066664f
C1488 diff_gen_0.delay_unit_2_6.in_2.t12 VSS 0.021266f
C1489 diff_gen_0.delay_unit_2_6.in_2.n4 VSS 0.046454f
C1490 diff_gen_0.delay_unit_2_6.in_2.n5 VSS 0.014821f
C1491 diff_gen_0.delay_unit_2_6.in_2.n6 VSS 0.22891f
C1492 diff_gen_0.delay_unit_2_6.in_2.t1 VSS 0.165681f
C1493 diff_gen_0.delay_unit_2_6.in_2.t0 VSS 0.051203f
C1494 diff_gen_0.delay_unit_2_6.in_2.n7 VSS 0.452839f
C1495 diff_gen_0.delay_unit_2_6.in_2.n8 VSS 0.285821f
C1496 diff_gen_0.delay_unit_2_6.in_2.t7 VSS 0.043739f
C1497 diff_gen_0.delay_unit_2_6.in_2.t5 VSS 0.043739f
C1498 diff_gen_0.delay_unit_2_6.in_2.n9 VSS 0.093535f
C1499 diff_gen_0.delay_unit_2_6.in_2.t3 VSS 0.01458f
C1500 diff_gen_0.delay_unit_2_6.in_2.t4 VSS 0.01458f
C1501 diff_gen_0.delay_unit_2_6.in_2.n10 VSS 0.031652f
C1502 diff_gen_0.delay_unit_2_6.in_2.n11 VSS 0.376142f
C1503 diff_gen_0.delay_unit_2_6.in_2.t6 VSS 0.165681f
C1504 diff_gen_0.delay_unit_2_6.in_2.t2 VSS 0.051203f
C1505 diff_gen_0.delay_unit_2_6.in_2.n12 VSS 0.398173f
C1506 diff_gen_0.delay_unit_2_6.in_2.n13 VSS 0.085944f
C1507 diff_gen_0.delay_unit_2_5.out_2 VSS 0.028637f
C1508 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1509 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1510 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.087567f
C1511 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.039891f
C1512 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1513 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C1514 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C1515 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.095888f
C1516 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.041221f
C1517 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C1518 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.108538f
C1519 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.081767f
C1520 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.090596f
C1521 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C1522 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C1523 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C1524 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C1525 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1526 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C1527 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.087824f
C1528 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.040008f
C1529 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C1530 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C1531 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.202807f
C1532 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.096169f
C1533 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.041341f
C1534 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C1535 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.082007f
C1536 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.090862f
C1537 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C1538 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C1539 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.107599f
C1540 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C1541 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.054421f
C1542 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C1543 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C1544 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
C1545 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t19 VSS 0.039259f
C1546 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t11 VSS 0.012524f
C1547 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n0 VSS 0.027535f
C1548 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t13 VSS 0.039259f
C1549 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t16 VSS 0.012524f
C1550 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1551 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1552 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t17 VSS 0.039259f
C1553 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t18 VSS 0.012524f
C1554 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n3 VSS 0.027535f
C1555 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t10 VSS 0.039259f
C1556 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t12 VSS 0.012524f
C1557 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1558 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1559 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1560 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t1 VSS 0.09757f
C1561 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t0 VSS 0.030153f
C1562 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1563 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t8 VSS 0.046129f
C1564 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t14 VSS 0.046129f
C1565 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1566 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t9 VSS 0.046129f
C1567 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t15 VSS 0.046129f
C1568 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1569 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1570 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t5 VSS 0.025758f
C1571 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t2 VSS 0.025758f
C1572 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1573 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t6 VSS 0.008586f
C1574 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t3 VSS 0.008586f
C1575 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1576 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1577 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t7 VSS 0.09757f
C1578 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.t4 VSS 0.030153f
C1579 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1580 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_2.n15 VSS 0.122976f
C1581 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t13 VSS 0.059856f
C1582 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t15 VSS 0.019094f
C1583 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n0 VSS 0.041709f
C1584 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t17 VSS 0.059856f
C1585 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t10 VSS 0.019094f
C1586 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n1 VSS 0.04198f
C1587 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n2 VSS 0.013454f
C1588 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t14 VSS 0.059856f
C1589 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t16 VSS 0.019094f
C1590 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n3 VSS 0.04198f
C1591 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t8 VSS 0.059856f
C1592 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t11 VSS 0.019094f
C1593 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n4 VSS 0.041709f
C1594 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n5 VSS 0.013307f
C1595 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n6 VSS 0.351208f
C1596 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t1 VSS 0.047903f
C1597 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t0 VSS 0.144997f
C1598 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n7 VSS 0.368007f
C1599 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n8 VSS 0.191794f
C1600 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t4 VSS 0.013091f
C1601 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t2 VSS 0.013091f
C1602 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n9 VSS 0.030662f
C1603 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t7 VSS 0.039272f
C1604 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t5 VSS 0.039272f
C1605 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n10 VSS 0.080004f
C1606 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n11 VSS 0.332866f
C1607 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t19 VSS 0.061472f
C1608 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t12 VSS 0.061472f
C1609 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n12 VSS 0.069399f
C1610 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t18 VSS 0.061472f
C1611 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t9 VSS 0.061472f
C1612 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n13 VSS 0.069022f
C1613 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n14 VSS 0.63019f
C1614 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t3 VSS 0.045973f
C1615 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n15 VSS 0.158781f
C1616 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.t6 VSS 0.144997f
C1617 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n16 VSS 0.240639f
C1618 vernier_delay_line_0.saff_delay_unit_4/delay_unit_2_0.in_1.n17 VSS 0.180864f
C1619 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.d VSS 0.696698f
C1620 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t8 VSS 0.059856f
C1621 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t11 VSS 0.019094f
C1622 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n0 VSS 0.041709f
C1623 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t13 VSS 0.059856f
C1624 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t16 VSS 0.019094f
C1625 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n1 VSS 0.04198f
C1626 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n2 VSS 0.013454f
C1627 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t19 VSS 0.059856f
C1628 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t10 VSS 0.019094f
C1629 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n3 VSS 0.04198f
C1630 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t15 VSS 0.059856f
C1631 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t18 VSS 0.019094f
C1632 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n4 VSS 0.041709f
C1633 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n5 VSS 0.013307f
C1634 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n6 VSS 0.351208f
C1635 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t0 VSS 0.047903f
C1636 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t1 VSS 0.144997f
C1637 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n7 VSS 0.368007f
C1638 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n8 VSS 0.191794f
C1639 vernier_delay_line_0.delay_unit_2_0.in_1 VSS 0.184027f
C1640 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t3 VSS 0.013091f
C1641 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t2 VSS 0.013091f
C1642 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n9 VSS 0.030662f
C1643 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t5 VSS 0.039272f
C1644 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t7 VSS 0.039272f
C1645 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n10 VSS 0.080004f
C1646 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n11 VSS 0.332866f
C1647 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t12 VSS 0.061472f
C1648 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t17 VSS 0.061472f
C1649 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n12 VSS 0.069399f
C1650 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t9 VSS 0.061472f
C1651 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t14 VSS 0.061472f
C1652 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n13 VSS 0.069022f
C1653 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n14 VSS 0.63019f
C1654 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t4 VSS 0.045973f
C1655 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n15 VSS 0.158781f
C1656 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.t6 VSS 0.144997f
C1657 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n16 VSS 0.240639f
C1658 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.d.n17 VSS 0.180864f
C1659 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_1 VSS 0.271416f
C1660 a_1082_2192.t7 VSS 0.024913f
C1661 a_1082_2192.t6 VSS 0.024913f
C1662 a_1082_2192.t5 VSS 0.024913f
C1663 a_1082_2192.n0 VSS 0.060272f
C1664 a_1082_2192.t3 VSS 0.024913f
C1665 a_1082_2192.t12 VSS 0.024913f
C1666 a_1082_2192.n1 VSS 0.060114f
C1667 a_1082_2192.t9 VSS 0.024913f
C1668 a_1082_2192.t11 VSS 0.024913f
C1669 a_1082_2192.n2 VSS 0.060114f
C1670 a_1082_2192.t1 VSS 0.024913f
C1671 a_1082_2192.t10 VSS 0.024913f
C1672 a_1082_2192.n3 VSS 0.060114f
C1673 a_1082_2192.t0 VSS 0.097139f
C1674 a_1082_2192.n4 VSS 0.369186f
C1675 a_1082_2192.n5 VSS 0.182473f
C1676 a_1082_2192.n6 VSS 0.22019f
C1677 a_1082_2192.t4 VSS 0.024913f
C1678 a_1082_2192.t2 VSS 0.024913f
C1679 a_1082_2192.n7 VSS 0.052659f
C1680 a_1082_2192.n8 VSS 0.140942f
C1681 a_1082_2192.n9 VSS 0.340434f
C1682 a_1082_2192.n10 VSS 0.057409f
C1683 a_1082_2192.t8 VSS 0.024913f
C1684 a_15038_2192.t2 VSS 0.059028f
C1685 a_15038_2192.t0 VSS 0.059028f
C1686 a_15038_2192.t1 VSS 0.059028f
C1687 a_15038_2192.n0 VSS 0.139449f
C1688 a_15038_2192.t5 VSS 0.059028f
C1689 a_15038_2192.t3 VSS 0.059028f
C1690 a_15038_2192.n1 VSS 0.258102f
C1691 a_15038_2192.n2 VSS 1.11221f
C1692 a_15038_2192.n3 VSS 0.136068f
C1693 a_15038_2192.t4 VSS 0.059028f
C1694 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t17 VSS 0.039259f
C1695 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t9 VSS 0.012524f
C1696 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n0 VSS 0.027534f
C1697 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t19 VSS 0.039259f
C1698 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t13 VSS 0.012524f
C1699 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1700 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1701 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t15 VSS 0.039259f
C1702 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t18 VSS 0.012524f
C1703 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n3 VSS 0.027534f
C1704 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t11 VSS 0.039259f
C1705 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t14 VSS 0.012524f
C1706 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1707 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1708 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1709 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t7 VSS 0.09757f
C1710 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t6 VSS 0.030153f
C1711 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1712 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t8 VSS 0.046129f
C1713 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t12 VSS 0.046129f
C1714 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1715 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t10 VSS 0.046129f
C1716 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t16 VSS 0.046129f
C1717 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1718 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1719 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t5 VSS 0.025758f
C1720 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t4 VSS 0.025758f
C1721 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1722 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t2 VSS 0.008586f
C1723 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t1 VSS 0.008586f
C1724 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1725 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1726 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t3 VSS 0.09757f
C1727 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.t0 VSS 0.030153f
C1728 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1729 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n15 VSS 0.050613f
C1730 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_2.n16 VSS 0.122976f
C1731 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C1732 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C1733 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.087567f
C1734 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.039891f
C1735 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C1736 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C1737 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.201734f
C1738 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.095888f
C1739 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.041221f
C1740 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C1741 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.108538f
C1742 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.081767f
C1743 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.090596f
C1744 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C1745 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.054262f
C1746 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C1747 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C1748 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C1749 diff_gen_0.delay_unit_2_5.in_1.t9 VSS 0.086195f
C1750 diff_gen_0.delay_unit_2_5.in_1.t12 VSS 0.027496f
C1751 diff_gen_0.delay_unit_2_5.in_1.n0 VSS 0.060063f
C1752 diff_gen_0.delay_unit_2_5.in_1.t8 VSS 0.086195f
C1753 diff_gen_0.delay_unit_2_5.in_1.t11 VSS 0.027496f
C1754 diff_gen_0.delay_unit_2_5.in_1.n1 VSS 0.060453f
C1755 diff_gen_0.delay_unit_2_5.in_1.n2 VSS 0.019374f
C1756 diff_gen_0.delay_unit_2_5.in_1.t15 VSS 0.086195f
C1757 diff_gen_0.delay_unit_2_5.in_1.t10 VSS 0.027496f
C1758 diff_gen_0.delay_unit_2_5.in_1.n3 VSS 0.060453f
C1759 diff_gen_0.delay_unit_2_5.in_1.t13 VSS 0.086195f
C1760 diff_gen_0.delay_unit_2_5.in_1.t14 VSS 0.027496f
C1761 diff_gen_0.delay_unit_2_5.in_1.n4 VSS 0.060063f
C1762 diff_gen_0.delay_unit_2_5.in_1.n5 VSS 0.019163f
C1763 diff_gen_0.delay_unit_2_5.in_1.n6 VSS 0.505752f
C1764 diff_gen_0.delay_unit_2_5.in_1.t3 VSS 0.068982f
C1765 diff_gen_0.delay_unit_2_5.in_1.t4 VSS 0.2088f
C1766 diff_gen_0.delay_unit_2_5.in_1.n7 VSS 0.529943f
C1767 diff_gen_0.delay_unit_2_5.in_1.n8 VSS 0.302399f
C1768 diff_gen_0.delay_unit_2_5.in_1.t2 VSS 0.018851f
C1769 diff_gen_0.delay_unit_2_5.in_1.t6 VSS 0.018851f
C1770 diff_gen_0.delay_unit_2_5.in_1.n9 VSS 0.044154f
C1771 diff_gen_0.delay_unit_2_5.in_1.t1 VSS 0.056553f
C1772 diff_gen_0.delay_unit_2_5.in_1.t0 VSS 0.056553f
C1773 diff_gen_0.delay_unit_2_5.in_1.n10 VSS 0.115209f
C1774 diff_gen_0.delay_unit_2_5.in_1.n11 VSS 0.479339f
C1775 diff_gen_0.delay_unit_2_5.in_1.t7 VSS 0.069002f
C1776 diff_gen_0.delay_unit_2_5.in_1.t5 VSS 0.2088f
C1777 diff_gen_0.delay_unit_2_5.in_1.n12 VSS 0.509237f
C1778 diff_gen_0.delay_unit_2_5.in_1.n13 VSS 0.26045f
C1779 diff_gen_0.delay_unit_2_4.out_1 VSS 0.212791f
C1780 a_3364_2192.t3 VSS 0.024913f
C1781 a_3364_2192.t4 VSS 0.024913f
C1782 a_3364_2192.t2 VSS 0.024913f
C1783 a_3364_2192.n0 VSS 0.057409f
C1784 a_3364_2192.t12 VSS 0.024913f
C1785 a_3364_2192.t9 VSS 0.024913f
C1786 a_3364_2192.n1 VSS 0.060114f
C1787 a_3364_2192.t7 VSS 0.024913f
C1788 a_3364_2192.t1 VSS 0.024913f
C1789 a_3364_2192.n2 VSS 0.060114f
C1790 a_3364_2192.t0 VSS 0.024913f
C1791 a_3364_2192.t10 VSS 0.024913f
C1792 a_3364_2192.n3 VSS 0.060114f
C1793 a_3364_2192.t8 VSS 0.097139f
C1794 a_3364_2192.n4 VSS 0.369186f
C1795 a_3364_2192.n5 VSS 0.182473f
C1796 a_3364_2192.n6 VSS 0.22019f
C1797 a_3364_2192.t5 VSS 0.024913f
C1798 a_3364_2192.t11 VSS 0.024913f
C1799 a_3364_2192.n7 VSS 0.052659f
C1800 a_3364_2192.n8 VSS 0.140942f
C1801 a_3364_2192.n9 VSS 0.340434f
C1802 a_3364_2192.n10 VSS 0.060272f
C1803 a_3364_2192.t6 VSS 0.024913f
C1804 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t13 VSS 0.059856f
C1805 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t16 VSS 0.019094f
C1806 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n0 VSS 0.041709f
C1807 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t18 VSS 0.059856f
C1808 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t9 VSS 0.019094f
C1809 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n1 VSS 0.04198f
C1810 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n2 VSS 0.013454f
C1811 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t19 VSS 0.059856f
C1812 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t10 VSS 0.019094f
C1813 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n3 VSS 0.04198f
C1814 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t11 VSS 0.059856f
C1815 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t15 VSS 0.019094f
C1816 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n4 VSS 0.041709f
C1817 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n5 VSS 0.013307f
C1818 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n6 VSS 0.351208f
C1819 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t0 VSS 0.047903f
C1820 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t3 VSS 0.144997f
C1821 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n7 VSS 0.368007f
C1822 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t6 VSS 0.013091f
C1823 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t5 VSS 0.013091f
C1824 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n8 VSS 0.030662f
C1825 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t1 VSS 0.039272f
C1826 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t2 VSS 0.039272f
C1827 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n9 VSS 0.080004f
C1828 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n10 VSS 0.332866f
C1829 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t12 VSS 0.061472f
C1830 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t17 VSS 0.061472f
C1831 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n11 VSS 0.069399f
C1832 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t8 VSS 0.061472f
C1833 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t14 VSS 0.061472f
C1834 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n12 VSS 0.069022f
C1835 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n13 VSS 0.63019f
C1836 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t4 VSS 0.045973f
C1837 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n14 VSS 0.158781f
C1838 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.t7 VSS 0.144997f
C1839 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n15 VSS 0.240639f
C1840 vernier_delay_line_0.saff_delay_unit_2/delay_unit_2_0.in_1.n16 VSS 0.180864f
C1841 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t10 VSS 0.039259f
C1842 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t13 VSS 0.012524f
C1843 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n0 VSS 0.027535f
C1844 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t16 VSS 0.039259f
C1845 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t19 VSS 0.012524f
C1846 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1847 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1848 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t8 VSS 0.039259f
C1849 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t11 VSS 0.012524f
C1850 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n3 VSS 0.027535f
C1851 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t14 VSS 0.039259f
C1852 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t17 VSS 0.012524f
C1853 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1854 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1855 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1856 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t0 VSS 0.09757f
C1857 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t1 VSS 0.030153f
C1858 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1859 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t9 VSS 0.046129f
C1860 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t15 VSS 0.046129f
C1861 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1862 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t12 VSS 0.046129f
C1863 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t18 VSS 0.046129f
C1864 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1865 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1866 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t3 VSS 0.025758f
C1867 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t5 VSS 0.025758f
C1868 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1869 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t4 VSS 0.008586f
C1870 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t2 VSS 0.008586f
C1871 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1872 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1873 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t7 VSS 0.09757f
C1874 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.t6 VSS 0.030153f
C1875 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1876 vernier_delay_line_0.saff_delay_unit_5/delay_unit_2_0.in_2.n15 VSS 0.122976f
C1877 a_5910_2192.t5 VSS 0.059028f
C1878 a_5910_2192.t0 VSS 0.059028f
C1879 a_5910_2192.t1 VSS 0.059028f
C1880 a_5910_2192.n0 VSS 0.139449f
C1881 a_5910_2192.t2 VSS 0.059028f
C1882 a_5910_2192.t3 VSS 0.059028f
C1883 a_5910_2192.n1 VSS 0.136068f
C1884 a_5910_2192.n2 VSS 1.11221f
C1885 a_5910_2192.n3 VSS 0.258102f
C1886 a_5910_2192.t4 VSS 0.059028f
C1887 a_5646_2192.t1 VSS 0.024913f
C1888 a_5646_2192.t0 VSS 0.024913f
C1889 a_5646_2192.t3 VSS 0.024913f
C1890 a_5646_2192.n0 VSS 0.060272f
C1891 a_5646_2192.t10 VSS 0.024913f
C1892 a_5646_2192.t6 VSS 0.024913f
C1893 a_5646_2192.n1 VSS 0.060114f
C1894 a_5646_2192.t7 VSS 0.024913f
C1895 a_5646_2192.t8 VSS 0.024913f
C1896 a_5646_2192.n2 VSS 0.060114f
C1897 a_5646_2192.t9 VSS 0.024913f
C1898 a_5646_2192.t5 VSS 0.024913f
C1899 a_5646_2192.n3 VSS 0.060114f
C1900 a_5646_2192.t12 VSS 0.097139f
C1901 a_5646_2192.n4 VSS 0.369186f
C1902 a_5646_2192.n5 VSS 0.182473f
C1903 a_5646_2192.n6 VSS 0.22019f
C1904 a_5646_2192.t2 VSS 0.024913f
C1905 a_5646_2192.t11 VSS 0.024913f
C1906 a_5646_2192.n7 VSS 0.052659f
C1907 a_5646_2192.n8 VSS 0.140942f
C1908 a_5646_2192.n9 VSS 0.340434f
C1909 a_5646_2192.n10 VSS 0.057409f
C1910 a_5646_2192.t4 VSS 0.024913f
C1911 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t13 VSS 0.039259f
C1912 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t15 VSS 0.012524f
C1913 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n0 VSS 0.027534f
C1914 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t9 VSS 0.039259f
C1915 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t11 VSS 0.012524f
C1916 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n1 VSS 0.027357f
C1917 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n2 VSS 0.008823f
C1918 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t14 VSS 0.039259f
C1919 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t17 VSS 0.012524f
C1920 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n3 VSS 0.027534f
C1921 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t16 VSS 0.039259f
C1922 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t19 VSS 0.012524f
C1923 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n4 VSS 0.027357f
C1924 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n5 VSS 0.008728f
C1925 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n6 VSS 0.134806f
C1926 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t6 VSS 0.09757f
C1927 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t5 VSS 0.030153f
C1928 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n7 VSS 0.266679f
C1929 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t10 VSS 0.046129f
C1930 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t8 VSS 0.046129f
C1931 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n8 VSS 0.054044f
C1932 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t18 VSS 0.046129f
C1933 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t12 VSS 0.046129f
C1934 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n9 VSS 0.0538f
C1935 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n10 VSS 0.493085f
C1936 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t1 VSS 0.025758f
C1937 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t2 VSS 0.025758f
C1938 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n11 VSS 0.055083f
C1939 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t3 VSS 0.008586f
C1940 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t7 VSS 0.008586f
C1941 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n12 VSS 0.01864f
C1942 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n13 VSS 0.221512f
C1943 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t4 VSS 0.09757f
C1944 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.t0 VSS 0.030153f
C1945 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n14 VSS 0.234486f
C1946 vernier_delay_line_0.saff_delay_unit_3/delay_unit_2_0.in_2.n15 VSS 0.122976f
C1947 vernier_delay_line_0.start_neg.t12 VSS 0.061832f
C1948 vernier_delay_line_0.start_neg.t14 VSS 0.019725f
C1949 vernier_delay_line_0.start_neg.n0 VSS 0.043367f
C1950 vernier_delay_line_0.start_neg.t8 VSS 0.061832f
C1951 vernier_delay_line_0.start_neg.t10 VSS 0.019725f
C1952 vernier_delay_line_0.start_neg.n1 VSS 0.043087f
C1953 vernier_delay_line_0.start_neg.n2 VSS 0.013896f
C1954 vernier_delay_line_0.start_neg.t11 VSS 0.061832f
C1955 vernier_delay_line_0.start_neg.t13 VSS 0.019725f
C1956 vernier_delay_line_0.start_neg.n3 VSS 0.043367f
C1957 vernier_delay_line_0.start_neg.t15 VSS 0.061832f
C1958 vernier_delay_line_0.start_neg.t9 VSS 0.019725f
C1959 vernier_delay_line_0.start_neg.n4 VSS 0.043087f
C1960 vernier_delay_line_0.start_neg.n5 VSS 0.013747f
C1961 vernier_delay_line_0.start_neg.n6 VSS 0.186471f
C1962 vernier_delay_line_0.start_neg.t6 VSS 0.153672f
C1963 vernier_delay_line_0.start_neg.t7 VSS 0.047491f
C1964 vernier_delay_line_0.start_neg.n7 VSS 0.420016f
C1965 vernier_delay_line_0.start_neg.t5 VSS 0.040569f
C1966 vernier_delay_line_0.start_neg.t3 VSS 0.040569f
C1967 vernier_delay_line_0.start_neg.n8 VSS 0.086755f
C1968 vernier_delay_line_0.start_neg.t0 VSS 0.013523f
C1969 vernier_delay_line_0.start_neg.t1 VSS 0.013523f
C1970 vernier_delay_line_0.start_neg.n9 VSS 0.029358f
C1971 vernier_delay_line_0.start_neg.n10 VSS 0.348878f
C1972 vernier_delay_line_0.start_neg.t4 VSS 0.153672f
C1973 vernier_delay_line_0.start_neg.t2 VSS 0.047491f
C1974 vernier_delay_line_0.start_neg.n11 VSS 0.369312f
C1975 vernier_delay_line_0.start_neg.n12 VSS 0.079715f
C1976 diff_gen_0.delay_unit_2_4.in_1.t13 VSS 0.086195f
C1977 diff_gen_0.delay_unit_2_4.in_1.t15 VSS 0.027496f
C1978 diff_gen_0.delay_unit_2_4.in_1.n0 VSS 0.060063f
C1979 diff_gen_0.delay_unit_2_4.in_1.t9 VSS 0.086195f
C1980 diff_gen_0.delay_unit_2_4.in_1.t11 VSS 0.027496f
C1981 diff_gen_0.delay_unit_2_4.in_1.n1 VSS 0.060453f
C1982 diff_gen_0.delay_unit_2_4.in_1.n2 VSS 0.019374f
C1983 diff_gen_0.delay_unit_2_4.in_1.t14 VSS 0.086195f
C1984 diff_gen_0.delay_unit_2_4.in_1.t8 VSS 0.027496f
C1985 diff_gen_0.delay_unit_2_4.in_1.n3 VSS 0.060453f
C1986 diff_gen_0.delay_unit_2_4.in_1.t10 VSS 0.086195f
C1987 diff_gen_0.delay_unit_2_4.in_1.t12 VSS 0.027496f
C1988 diff_gen_0.delay_unit_2_4.in_1.n4 VSS 0.060063f
C1989 diff_gen_0.delay_unit_2_4.in_1.n5 VSS 0.019163f
C1990 diff_gen_0.delay_unit_2_4.in_1.n6 VSS 0.505752f
C1991 diff_gen_0.delay_unit_2_4.in_1.t0 VSS 0.068982f
C1992 diff_gen_0.delay_unit_2_4.in_1.t7 VSS 0.2088f
C1993 diff_gen_0.delay_unit_2_4.in_1.n7 VSS 0.529943f
C1994 diff_gen_0.delay_unit_2_4.in_1.n8 VSS 0.27619f
C1995 diff_gen_0.delay_unit_2_4.in_1.t3 VSS 0.018851f
C1996 diff_gen_0.delay_unit_2_4.in_1.t1 VSS 0.018851f
C1997 diff_gen_0.delay_unit_2_4.in_1.n9 VSS 0.044154f
C1998 diff_gen_0.delay_unit_2_4.in_1.t6 VSS 0.056553f
C1999 diff_gen_0.delay_unit_2_4.in_1.t4 VSS 0.056553f
C2000 diff_gen_0.delay_unit_2_4.in_1.n10 VSS 0.115209f
C2001 diff_gen_0.delay_unit_2_4.in_1.n11 VSS 0.479339f
C2002 diff_gen_0.delay_unit_2_4.in_1.t2 VSS 0.069002f
C2003 diff_gen_0.delay_unit_2_4.in_1.t5 VSS 0.2088f
C2004 diff_gen_0.delay_unit_2_4.in_1.n12 VSS 0.509237f
C2005 diff_gen_0.delay_unit_2_4.in_1.n13 VSS 0.26045f
C2006 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t13 VSS 0.039259f
C2007 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t15 VSS 0.012524f
C2008 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n0 VSS 0.027535f
C2009 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t17 VSS 0.039259f
C2010 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t8 VSS 0.012524f
C2011 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n1 VSS 0.027357f
C2012 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n2 VSS 0.008823f
C2013 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t10 VSS 0.039259f
C2014 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t14 VSS 0.012524f
C2015 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n3 VSS 0.027535f
C2016 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t19 VSS 0.039259f
C2017 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t9 VSS 0.012524f
C2018 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n4 VSS 0.027357f
C2019 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n5 VSS 0.008728f
C2020 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n6 VSS 0.134806f
C2021 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t1 VSS 0.09757f
C2022 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t0 VSS 0.030153f
C2023 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n7 VSS 0.266679f
C2024 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t11 VSS 0.046129f
C2025 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t16 VSS 0.046129f
C2026 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n8 VSS 0.054044f
C2027 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t18 VSS 0.046129f
C2028 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t12 VSS 0.046129f
C2029 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n9 VSS 0.0538f
C2030 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n10 VSS 0.493085f
C2031 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t2 VSS 0.025758f
C2032 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t6 VSS 0.025758f
C2033 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n11 VSS 0.055083f
C2034 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t4 VSS 0.008586f
C2035 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t3 VSS 0.008586f
C2036 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n12 VSS 0.01864f
C2037 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n13 VSS 0.221512f
C2038 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t5 VSS 0.09757f
C2039 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.t7 VSS 0.030153f
C2040 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n14 VSS 0.234486f
C2041 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_2.n15 VSS 0.122976f
C2042 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t14 VSS 0.059856f
C2043 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t19 VSS 0.019094f
C2044 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n0 VSS 0.041709f
C2045 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t9 VSS 0.059856f
C2046 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t11 VSS 0.019094f
C2047 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n1 VSS 0.04198f
C2048 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n2 VSS 0.013454f
C2049 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t12 VSS 0.059856f
C2050 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t17 VSS 0.019094f
C2051 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n3 VSS 0.04198f
C2052 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t15 VSS 0.059856f
C2053 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t8 VSS 0.019094f
C2054 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n4 VSS 0.041709f
C2055 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n5 VSS 0.013307f
C2056 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n6 VSS 0.351208f
C2057 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t7 VSS 0.047903f
C2058 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t6 VSS 0.144997f
C2059 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n7 VSS 0.368007f
C2060 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t1 VSS 0.013091f
C2061 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t4 VSS 0.013091f
C2062 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n8 VSS 0.030662f
C2063 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t5 VSS 0.039272f
C2064 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t0 VSS 0.039272f
C2065 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n9 VSS 0.080004f
C2066 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n10 VSS 0.332866f
C2067 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t13 VSS 0.061472f
C2068 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t18 VSS 0.061472f
C2069 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n11 VSS 0.069399f
C2070 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t10 VSS 0.061472f
C2071 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t16 VSS 0.061472f
C2072 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n12 VSS 0.069022f
C2073 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n13 VSS 0.63019f
C2074 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t2 VSS 0.045973f
C2075 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n14 VSS 0.158781f
C2076 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.t3 VSS 0.144997f
C2077 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n15 VSS 0.240639f
C2078 vernier_delay_line_0.saff_delay_unit_6/delay_unit_2_0.in_1.n16 VSS 0.180864f
C2079 diff_gen_0.delay_unit_2_1.in_1.t10 VSS 0.086195f
C2080 diff_gen_0.delay_unit_2_1.in_1.t13 VSS 0.027496f
C2081 diff_gen_0.delay_unit_2_1.in_1.n0 VSS 0.060063f
C2082 diff_gen_0.delay_unit_2_1.in_1.t15 VSS 0.086195f
C2083 diff_gen_0.delay_unit_2_1.in_1.t8 VSS 0.027496f
C2084 diff_gen_0.delay_unit_2_1.in_1.n1 VSS 0.060453f
C2085 diff_gen_0.delay_unit_2_1.in_1.n2 VSS 0.019374f
C2086 diff_gen_0.delay_unit_2_1.in_1.t11 VSS 0.086195f
C2087 diff_gen_0.delay_unit_2_1.in_1.t14 VSS 0.027496f
C2088 diff_gen_0.delay_unit_2_1.in_1.n3 VSS 0.060453f
C2089 diff_gen_0.delay_unit_2_1.in_1.t9 VSS 0.086195f
C2090 diff_gen_0.delay_unit_2_1.in_1.t12 VSS 0.027496f
C2091 diff_gen_0.delay_unit_2_1.in_1.n4 VSS 0.060063f
C2092 diff_gen_0.delay_unit_2_1.in_1.n5 VSS 0.019163f
C2093 diff_gen_0.delay_unit_2_1.in_1.n6 VSS 0.505752f
C2094 diff_gen_0.delay_unit_2_1.in_1.t0 VSS 0.068982f
C2095 diff_gen_0.delay_unit_2_1.in_1.t1 VSS 0.2088f
C2096 diff_gen_0.delay_unit_2_1.in_1.n7 VSS 0.529943f
C2097 diff_gen_0.delay_unit_2_1.in_1.n8 VSS 0.27619f
C2098 diff_gen_0.delay_unit_2_1.in_1.t2 VSS 0.018851f
C2099 diff_gen_0.delay_unit_2_1.in_1.t3 VSS 0.018851f
C2100 diff_gen_0.delay_unit_2_1.in_1.n9 VSS 0.044154f
C2101 diff_gen_0.delay_unit_2_1.in_1.t5 VSS 0.056553f
C2102 diff_gen_0.delay_unit_2_1.in_1.t6 VSS 0.056553f
C2103 diff_gen_0.delay_unit_2_1.in_1.n10 VSS 0.115209f
C2104 diff_gen_0.delay_unit_2_1.in_1.n11 VSS 0.479339f
C2105 diff_gen_0.delay_unit_2_1.in_1.t4 VSS 0.069002f
C2106 diff_gen_0.delay_unit_2_1.in_1.t7 VSS 0.2088f
C2107 diff_gen_0.delay_unit_2_1.in_1.n12 VSS 0.509237f
C2108 diff_gen_0.delay_unit_2_1.in_1.n13 VSS 0.26045f
C2109 diff_gen_0.delay_unit_2_1.in_2.t10 VSS 0.066664f
C2110 diff_gen_0.delay_unit_2_1.in_2.t12 VSS 0.021266f
C2111 diff_gen_0.delay_unit_2_1.in_2.n0 VSS 0.046756f
C2112 diff_gen_0.delay_unit_2_1.in_2.t15 VSS 0.066664f
C2113 diff_gen_0.delay_unit_2_1.in_2.t9 VSS 0.021266f
C2114 diff_gen_0.delay_unit_2_1.in_2.n1 VSS 0.046454f
C2115 diff_gen_0.delay_unit_2_1.in_2.n2 VSS 0.014982f
C2116 diff_gen_0.delay_unit_2_1.in_2.t11 VSS 0.066664f
C2117 diff_gen_0.delay_unit_2_1.in_2.t13 VSS 0.021266f
C2118 diff_gen_0.delay_unit_2_1.in_2.n3 VSS 0.046756f
C2119 diff_gen_0.delay_unit_2_1.in_2.t14 VSS 0.066664f
C2120 diff_gen_0.delay_unit_2_1.in_2.t8 VSS 0.021266f
C2121 diff_gen_0.delay_unit_2_1.in_2.n4 VSS 0.046454f
C2122 diff_gen_0.delay_unit_2_1.in_2.n5 VSS 0.014821f
C2123 diff_gen_0.delay_unit_2_1.in_2.n6 VSS 0.22891f
C2124 diff_gen_0.delay_unit_2_1.in_2.t7 VSS 0.165681f
C2125 diff_gen_0.delay_unit_2_1.in_2.t0 VSS 0.051203f
C2126 diff_gen_0.delay_unit_2_1.in_2.n7 VSS 0.452839f
C2127 diff_gen_0.delay_unit_2_1.in_2.n8 VSS 0.285821f
C2128 diff_gen_0.delay_unit_2_1.in_2.t4 VSS 0.043739f
C2129 diff_gen_0.delay_unit_2_1.in_2.t5 VSS 0.043739f
C2130 diff_gen_0.delay_unit_2_1.in_2.n9 VSS 0.093535f
C2131 diff_gen_0.delay_unit_2_1.in_2.t3 VSS 0.01458f
C2132 diff_gen_0.delay_unit_2_1.in_2.t1 VSS 0.01458f
C2133 diff_gen_0.delay_unit_2_1.in_2.n10 VSS 0.031652f
C2134 diff_gen_0.delay_unit_2_1.in_2.n11 VSS 0.376142f
C2135 diff_gen_0.delay_unit_2_1.in_2.t6 VSS 0.165681f
C2136 diff_gen_0.delay_unit_2_1.in_2.t2 VSS 0.051203f
C2137 diff_gen_0.delay_unit_2_1.in_2.n12 VSS 0.398173f
C2138 diff_gen_0.delay_unit_2_1.in_2.n13 VSS 0.085944f
C2139 diff_gen_0.delay_unit_2_0.out_2 VSS 0.028637f
C2140 a_n6458_3464.t6 VSS 0.228995f
C2141 a_n6458_3464.t35 VSS 0.093349f
C2142 a_n6458_3464.t38 VSS 0.030133f
C2143 a_n6458_3464.n0 VSS 0.086421f
C2144 a_n6458_3464.t28 VSS 0.093349f
C2145 a_n6458_3464.t29 VSS 0.030133f
C2146 a_n6458_3464.n1 VSS 0.088816f
C2147 a_n6458_3464.t11 VSS 0.093349f
C2148 a_n6458_3464.t14 VSS 0.030133f
C2149 a_n6458_3464.n2 VSS 0.088354f
C2150 a_n6458_3464.n3 VSS 0.389976f
C2151 a_n6458_3464.t33 VSS 0.093349f
C2152 a_n6458_3464.t36 VSS 0.030133f
C2153 a_n6458_3464.n4 VSS 0.088354f
C2154 a_n6458_3464.n5 VSS 0.217864f
C2155 a_n6458_3464.t23 VSS 0.093349f
C2156 a_n6458_3464.t25 VSS 0.030133f
C2157 a_n6458_3464.n6 VSS 0.088354f
C2158 a_n6458_3464.n7 VSS 0.217864f
C2159 a_n6458_3464.t15 VSS 0.093349f
C2160 a_n6458_3464.t18 VSS 0.030133f
C2161 a_n6458_3464.n8 VSS 0.088354f
C2162 a_n6458_3464.n9 VSS 0.217864f
C2163 a_n6458_3464.t37 VSS 0.093349f
C2164 a_n6458_3464.t39 VSS 0.030133f
C2165 a_n6458_3464.n10 VSS 0.088354f
C2166 a_n6458_3464.n11 VSS 0.217864f
C2167 a_n6458_3464.t26 VSS 0.093349f
C2168 a_n6458_3464.t27 VSS 0.030133f
C2169 a_n6458_3464.n12 VSS 0.088354f
C2170 a_n6458_3464.n13 VSS 0.217864f
C2171 a_n6458_3464.t19 VSS 0.093349f
C2172 a_n6458_3464.t22 VSS 0.030133f
C2173 a_n6458_3464.n14 VSS 0.088354f
C2174 a_n6458_3464.n15 VSS 0.217864f
C2175 a_n6458_3464.t8 VSS 0.093349f
C2176 a_n6458_3464.t9 VSS 0.030133f
C2177 a_n6458_3464.n16 VSS 0.088354f
C2178 a_n6458_3464.n17 VSS 0.217864f
C2179 a_n6458_3464.t30 VSS 0.093349f
C2180 a_n6458_3464.t31 VSS 0.030133f
C2181 a_n6458_3464.n18 VSS 0.088354f
C2182 a_n6458_3464.n19 VSS 0.217864f
C2183 a_n6458_3464.t17 VSS 0.093349f
C2184 a_n6458_3464.t20 VSS 0.030133f
C2185 a_n6458_3464.n20 VSS 0.088354f
C2186 a_n6458_3464.n21 VSS 0.217864f
C2187 a_n6458_3464.t10 VSS 0.093349f
C2188 a_n6458_3464.t12 VSS 0.030133f
C2189 a_n6458_3464.n22 VSS 0.088354f
C2190 a_n6458_3464.n23 VSS 0.217864f
C2191 a_n6458_3464.t32 VSS 0.093349f
C2192 a_n6458_3464.t34 VSS 0.030133f
C2193 a_n6458_3464.n24 VSS 0.088354f
C2194 a_n6458_3464.n25 VSS 0.217864f
C2195 a_n6458_3464.t21 VSS 0.093349f
C2196 a_n6458_3464.t24 VSS 0.030133f
C2197 a_n6458_3464.n26 VSS 0.088354f
C2198 a_n6458_3464.n27 VSS 0.217864f
C2199 a_n6458_3464.t13 VSS 0.093349f
C2200 a_n6458_3464.t16 VSS 0.030133f
C2201 a_n6458_3464.n28 VSS 0.088354f
C2202 a_n6458_3464.n29 VSS 0.289551f
C2203 a_n6458_3464.n30 VSS 0.109352f
C2204 a_n6458_3464.n31 VSS 0.42154f
C2205 a_n6458_3464.t1 VSS 0.071536f
C2206 a_n6458_3464.n32 VSS 0.133321f
C2207 a_n6458_3464.t4 VSS 0.231476f
C2208 a_n6458_3464.t3 VSS 0.071536f
C2209 a_n6458_3464.n33 VSS 0.529025f
C2210 a_n6458_3464.n34 VSS 0.22418f
C2211 a_n6458_3464.t5 VSS 0.231476f
C2212 a_n6458_3464.t0 VSS 0.071536f
C2213 a_n6458_3464.n35 VSS 0.538008f
C2214 a_n6458_3464.n36 VSS 0.22418f
C2215 a_n6458_3464.t2 VSS 0.071536f
C2216 a_n6458_3464.n37 VSS 0.529025f
C2217 a_n6458_3464.t7 VSS 0.231476f
C2218 vernier_delay_line_0.delay_unit_2_0.in_2 VSS 0.191438f
C2219 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t9 VSS 0.046129f
C2220 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t17 VSS 0.046129f
C2221 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n0 VSS 0.054044f
C2222 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t13 VSS 0.046129f
C2223 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t18 VSS 0.046129f
C2224 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n1 VSS 0.0538f
C2225 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n2 VSS 0.493085f
C2226 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.nd VSS 0.377104f
C2227 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t11 VSS 0.039259f
C2228 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t14 VSS 0.012524f
C2229 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n3 VSS 0.027534f
C2230 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t19 VSS 0.039259f
C2231 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t10 VSS 0.012524f
C2232 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n4 VSS 0.027357f
C2233 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n5 VSS 0.008823f
C2234 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t8 VSS 0.039259f
C2235 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t12 VSS 0.012524f
C2236 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n6 VSS 0.027534f
C2237 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t15 VSS 0.039259f
C2238 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t16 VSS 0.012524f
C2239 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n7 VSS 0.027357f
C2240 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n8 VSS 0.008728f
C2241 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n9 VSS 0.134806f
C2242 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t1 VSS 0.09757f
C2243 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t0 VSS 0.030153f
C2244 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n10 VSS 0.266679f
C2245 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n11 VSS 0.122976f
C2246 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t7 VSS 0.025758f
C2247 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t6 VSS 0.025758f
C2248 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n12 VSS 0.055083f
C2249 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t2 VSS 0.008586f
C2250 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t4 VSS 0.008586f
C2251 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n13 VSS 0.01864f
C2252 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n14 VSS 0.221512f
C2253 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t5 VSS 0.09757f
C2254 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.t3 VSS 0.030153f
C2255 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n15 VSS 0.234486f
C2256 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.nd.n16 VSS 0.050613f
C2257 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.out_2 VSS 0.082616f
C2258 start_buffer_0.start_delay.t6 VSS 0.1725f
C2259 start_buffer_0.start_delay.t2 VSS 0.05331f
C2260 start_buffer_0.start_delay.n0 VSS 0.400932f
C2261 start_buffer_0.start_delay.t5 VSS 0.1725f
C2262 start_buffer_0.start_delay.t1 VSS 0.05331f
C2263 start_buffer_0.start_delay.n1 VSS 0.394238f
C2264 start_buffer_0.start_delay.n2 VSS 0.167063f
C2265 start_buffer_0.start_delay.t4 VSS 0.170686f
C2266 start_buffer_0.start_delay.n3 VSS 0.310685f
C2267 start_buffer_0.start_delay.t0 VSS 0.05331f
C2268 start_buffer_0.start_delay.n4 VSS 0.09314f
C2269 start_buffer_0.start_delay.n5 VSS 0.131763f
C2270 start_buffer_0.start_delay.t8 VSS 0.069408f
C2271 start_buffer_0.start_delay.t10 VSS 0.022142f
C2272 start_buffer_0.start_delay.n6 VSS 0.04868f
C2273 start_buffer_0.start_delay.t12 VSS 0.069408f
C2274 start_buffer_0.start_delay.t15 VSS 0.022142f
C2275 start_buffer_0.start_delay.n7 VSS 0.048366f
C2276 start_buffer_0.start_delay.n8 VSS 0.015598f
C2277 start_buffer_0.start_delay.t11 VSS 0.069408f
C2278 start_buffer_0.start_delay.t13 VSS 0.022142f
C2279 start_buffer_0.start_delay.n9 VSS 0.04868f
C2280 start_buffer_0.start_delay.t14 VSS 0.069408f
C2281 start_buffer_0.start_delay.t9 VSS 0.022142f
C2282 start_buffer_0.start_delay.n10 VSS 0.048366f
C2283 start_buffer_0.start_delay.n11 VSS 0.015431f
C2284 start_buffer_0.start_delay.n12 VSS 0.188318f
C2285 start_buffer_0.start_delay.t7 VSS 0.1725f
C2286 start_buffer_0.start_delay.t3 VSS 0.05331f
C2287 start_buffer_0.start_delay.n13 VSS 0.471477f
C2288 start_buffer_0.start_buff.t11 VSS 0.07812f
C2289 start_buffer_0.start_buff.t14 VSS 0.024921f
C2290 start_buffer_0.start_buff.n0 VSS 0.054437f
C2291 start_buffer_0.start_buff.t21 VSS 0.07812f
C2292 start_buffer_0.start_buff.t12 VSS 0.024921f
C2293 start_buffer_0.start_buff.n1 VSS 0.05479f
C2294 start_buffer_0.start_buff.n2 VSS 0.017559f
C2295 start_buffer_0.start_buff.t17 VSS 0.07812f
C2296 start_buffer_0.start_buff.t18 VSS 0.024921f
C2297 start_buffer_0.start_buff.n3 VSS 0.05479f
C2298 start_buffer_0.start_buff.t10 VSS 0.07812f
C2299 start_buffer_0.start_buff.t13 VSS 0.024921f
C2300 start_buffer_0.start_buff.n4 VSS 0.054437f
C2301 start_buffer_0.start_buff.n5 VSS 0.017368f
C2302 start_buffer_0.start_buff.n6 VSS 0.458376f
C2303 start_buffer_0.start_buff.t8 VSS 0.06252f
C2304 start_buffer_0.start_buff.t9 VSS 0.189241f
C2305 start_buffer_0.start_buff.n7 VSS 0.480301f
C2306 start_buffer_0.start_buff.n8 VSS 0.250318f
C2307 start_buffer_0.start_buff.t5 VSS 0.189241f
C2308 start_buffer_0.start_buff.n9 VSS 0.429508f
C2309 start_buffer_0.start_buff.t15 VSS 0.078297f
C2310 start_buffer_0.start_buff.t16 VSS 0.025274f
C2311 start_buffer_0.start_buff.n10 VSS 0.072486f
C2312 start_buffer_0.start_buff.t22 VSS 0.078297f
C2313 start_buffer_0.start_buff.t23 VSS 0.025274f
C2314 start_buffer_0.start_buff.n11 VSS 0.074495f
C2315 start_buffer_0.start_buff.t19 VSS 0.078297f
C2316 start_buffer_0.start_buff.t20 VSS 0.025274f
C2317 start_buffer_0.start_buff.n12 VSS 0.074107f
C2318 start_buffer_0.start_buff.n13 VSS 0.387222f
C2319 start_buffer_0.start_buff.n14 VSS 0.091249f
C2320 start_buffer_0.start_buff.n15 VSS 0.089396f
C2321 start_buffer_0.start_buff.t0 VSS 0.060002f
C2322 start_buffer_0.start_buff.n16 VSS 0.10513f
C2323 start_buffer_0.start_buff.t4 VSS 0.194152f
C2324 start_buffer_0.start_buff.t3 VSS 0.060002f
C2325 start_buffer_0.start_buff.n17 VSS 0.451257f
C2326 start_buffer_0.start_buff.t7 VSS 0.194152f
C2327 start_buffer_0.start_buff.t2 VSS 0.060002f
C2328 start_buffer_0.start_buff.n18 VSS 0.443723f
C2329 start_buffer_0.start_buff.n19 VSS 0.188032f
C2330 start_buffer_0.start_buff.t6 VSS 0.194152f
C2331 start_buffer_0.start_buff.t1 VSS 0.060002f
C2332 start_buffer_0.start_buff.n20 VSS 0.443723f
C2333 start_buffer_0.start_buff.n21 VSS 0.113248f
C2334 diff_gen_0.delay_unit_2_3.in_2.t12 VSS 0.066664f
C2335 diff_gen_0.delay_unit_2_3.in_2.t14 VSS 0.021266f
C2336 diff_gen_0.delay_unit_2_3.in_2.n0 VSS 0.046756f
C2337 diff_gen_0.delay_unit_2_3.in_2.t8 VSS 0.066664f
C2338 diff_gen_0.delay_unit_2_3.in_2.t10 VSS 0.021266f
C2339 diff_gen_0.delay_unit_2_3.in_2.n1 VSS 0.046454f
C2340 diff_gen_0.delay_unit_2_3.in_2.n2 VSS 0.014982f
C2341 diff_gen_0.delay_unit_2_3.in_2.t13 VSS 0.066664f
C2342 diff_gen_0.delay_unit_2_3.in_2.t15 VSS 0.021266f
C2343 diff_gen_0.delay_unit_2_3.in_2.n3 VSS 0.046756f
C2344 diff_gen_0.delay_unit_2_3.in_2.t9 VSS 0.066664f
C2345 diff_gen_0.delay_unit_2_3.in_2.t11 VSS 0.021266f
C2346 diff_gen_0.delay_unit_2_3.in_2.n4 VSS 0.046454f
C2347 diff_gen_0.delay_unit_2_3.in_2.n5 VSS 0.014821f
C2348 diff_gen_0.delay_unit_2_3.in_2.n6 VSS 0.22891f
C2349 diff_gen_0.delay_unit_2_3.in_2.t7 VSS 0.165681f
C2350 diff_gen_0.delay_unit_2_3.in_2.t6 VSS 0.051203f
C2351 diff_gen_0.delay_unit_2_3.in_2.n7 VSS 0.452839f
C2352 diff_gen_0.delay_unit_2_3.in_2.n8 VSS 0.285821f
C2353 diff_gen_0.delay_unit_2_3.in_2.t3 VSS 0.043739f
C2354 diff_gen_0.delay_unit_2_3.in_2.t4 VSS 0.043739f
C2355 diff_gen_0.delay_unit_2_3.in_2.n9 VSS 0.093535f
C2356 diff_gen_0.delay_unit_2_3.in_2.t2 VSS 0.01458f
C2357 diff_gen_0.delay_unit_2_3.in_2.t0 VSS 0.01458f
C2358 diff_gen_0.delay_unit_2_3.in_2.n10 VSS 0.031652f
C2359 diff_gen_0.delay_unit_2_3.in_2.n11 VSS 0.376142f
C2360 diff_gen_0.delay_unit_2_3.in_2.t5 VSS 0.165681f
C2361 diff_gen_0.delay_unit_2_3.in_2.t1 VSS 0.051203f
C2362 diff_gen_0.delay_unit_2_3.in_2.n12 VSS 0.398173f
C2363 diff_gen_0.delay_unit_2_3.in_2.n13 VSS 0.085944f
C2364 diff_gen_0.delay_unit_2_2.out_2 VSS 0.028637f
C2365 diff_gen_0.delay_unit_2_2.in_1.t9 VSS 0.086195f
C2366 diff_gen_0.delay_unit_2_2.in_1.t12 VSS 0.027496f
C2367 diff_gen_0.delay_unit_2_2.in_1.n0 VSS 0.060063f
C2368 diff_gen_0.delay_unit_2_2.in_1.t15 VSS 0.086195f
C2369 diff_gen_0.delay_unit_2_2.in_1.t8 VSS 0.027496f
C2370 diff_gen_0.delay_unit_2_2.in_1.n1 VSS 0.060453f
C2371 diff_gen_0.delay_unit_2_2.in_1.n2 VSS 0.019374f
C2372 diff_gen_0.delay_unit_2_2.in_1.t11 VSS 0.086195f
C2373 diff_gen_0.delay_unit_2_2.in_1.t14 VSS 0.027496f
C2374 diff_gen_0.delay_unit_2_2.in_1.n3 VSS 0.060453f
C2375 diff_gen_0.delay_unit_2_2.in_1.t10 VSS 0.086195f
C2376 diff_gen_0.delay_unit_2_2.in_1.t13 VSS 0.027496f
C2377 diff_gen_0.delay_unit_2_2.in_1.n4 VSS 0.060063f
C2378 diff_gen_0.delay_unit_2_2.in_1.n5 VSS 0.019163f
C2379 diff_gen_0.delay_unit_2_2.in_1.n6 VSS 0.505752f
C2380 diff_gen_0.delay_unit_2_2.in_1.t6 VSS 0.068982f
C2381 diff_gen_0.delay_unit_2_2.in_1.t4 VSS 0.2088f
C2382 diff_gen_0.delay_unit_2_2.in_1.n7 VSS 0.529943f
C2383 diff_gen_0.delay_unit_2_2.in_1.n8 VSS 0.302399f
C2384 diff_gen_0.delay_unit_2_2.in_1.t5 VSS 0.018851f
C2385 diff_gen_0.delay_unit_2_2.in_1.t0 VSS 0.018851f
C2386 diff_gen_0.delay_unit_2_2.in_1.n9 VSS 0.044154f
C2387 diff_gen_0.delay_unit_2_2.in_1.t3 VSS 0.056553f
C2388 diff_gen_0.delay_unit_2_2.in_1.t2 VSS 0.056553f
C2389 diff_gen_0.delay_unit_2_2.in_1.n10 VSS 0.115209f
C2390 diff_gen_0.delay_unit_2_2.in_1.n11 VSS 0.479339f
C2391 diff_gen_0.delay_unit_2_2.in_1.t7 VSS 0.069002f
C2392 diff_gen_0.delay_unit_2_2.in_1.t1 VSS 0.2088f
C2393 diff_gen_0.delay_unit_2_2.in_1.n12 VSS 0.509237f
C2394 diff_gen_0.delay_unit_2_2.in_1.n13 VSS 0.26045f
C2395 diff_gen_0.delay_unit_2_1.out_1 VSS 0.212791f
C2396 a_12492_2192.t6 VSS 0.024913f
C2397 a_12492_2192.t7 VSS 0.024913f
C2398 a_12492_2192.t5 VSS 0.024913f
C2399 a_12492_2192.n0 VSS 0.060272f
C2400 a_12492_2192.t12 VSS 0.024913f
C2401 a_12492_2192.t3 VSS 0.024913f
C2402 a_12492_2192.n1 VSS 0.060114f
C2403 a_12492_2192.t2 VSS 0.024913f
C2404 a_12492_2192.t1 VSS 0.024913f
C2405 a_12492_2192.n2 VSS 0.060114f
C2406 a_12492_2192.t4 VSS 0.024913f
C2407 a_12492_2192.t0 VSS 0.024913f
C2408 a_12492_2192.n3 VSS 0.060114f
C2409 a_12492_2192.t10 VSS 0.097139f
C2410 a_12492_2192.n4 VSS 0.369186f
C2411 a_12492_2192.n5 VSS 0.182473f
C2412 a_12492_2192.n6 VSS 0.22019f
C2413 a_12492_2192.t8 VSS 0.024913f
C2414 a_12492_2192.t11 VSS 0.024913f
C2415 a_12492_2192.n7 VSS 0.052659f
C2416 a_12492_2192.n8 VSS 0.140942f
C2417 a_12492_2192.n9 VSS 0.340434f
C2418 a_12492_2192.n10 VSS 0.057409f
C2419 a_12492_2192.t9 VSS 0.024913f
C2420 stop_buffer_0.stop_strong VSS 0.454861f
C2421 vernier_delay_line_0.stop_strong.t79 VSS 0.093756f
C2422 vernier_delay_line_0.stop_strong.t75 VSS 0.093545f
C2423 vernier_delay_line_0.stop_strong.n0 VSS 0.403473f
C2424 vernier_delay_line_0.stop_strong.t72 VSS 0.072027f
C2425 vernier_delay_line_0.stop_strong.t38 VSS 0.072027f
C2426 vernier_delay_line_0.stop_strong.t43 VSS 0.072027f
C2427 vernier_delay_line_0.stop_strong.t59 VSS 0.072027f
C2428 vernier_delay_line_0.stop_strong.t80 VSS 0.079805f
C2429 vernier_delay_line_0.stop_strong.n1 VSS 0.070183f
C2430 vernier_delay_line_0.stop_strong.n2 VSS 0.04137f
C2431 vernier_delay_line_0.stop_strong.n3 VSS 0.04137f
C2432 vernier_delay_line_0.stop_strong.n4 VSS 0.062319f
C2433 vernier_delay_line_0.stop_strong.n5 VSS 0.937097f
C2434 vernier_delay_line_0.stop_strong.t21 VSS 0.181057f
C2435 vernier_delay_line_0.stop_strong.t16 VSS 0.055955f
C2436 vernier_delay_line_0.stop_strong.n6 VSS 0.420822f
C2437 vernier_delay_line_0.stop_strong.t9 VSS 0.181057f
C2438 vernier_delay_line_0.stop_strong.t14 VSS 0.055955f
C2439 vernier_delay_line_0.stop_strong.n7 VSS 0.413796f
C2440 vernier_delay_line_0.stop_strong.n8 VSS 0.17535f
C2441 vernier_delay_line_0.stop_strong.t3 VSS 0.181057f
C2442 vernier_delay_line_0.stop_strong.t28 VSS 0.055955f
C2443 vernier_delay_line_0.stop_strong.n9 VSS 0.413796f
C2444 vernier_delay_line_0.stop_strong.n10 VSS 0.11234f
C2445 vernier_delay_line_0.stop_strong.t18 VSS 0.181057f
C2446 vernier_delay_line_0.stop_strong.t20 VSS 0.055955f
C2447 vernier_delay_line_0.stop_strong.n11 VSS 0.413796f
C2448 vernier_delay_line_0.stop_strong.n12 VSS 0.11234f
C2449 vernier_delay_line_0.stop_strong.t6 VSS 0.181057f
C2450 vernier_delay_line_0.stop_strong.t8 VSS 0.055955f
C2451 vernier_delay_line_0.stop_strong.n13 VSS 0.413796f
C2452 vernier_delay_line_0.stop_strong.n14 VSS 0.11234f
C2453 vernier_delay_line_0.stop_strong.t15 VSS 0.181057f
C2454 vernier_delay_line_0.stop_strong.t2 VSS 0.055955f
C2455 vernier_delay_line_0.stop_strong.n15 VSS 0.413796f
C2456 vernier_delay_line_0.stop_strong.n16 VSS 0.11234f
C2457 vernier_delay_line_0.stop_strong.t0 VSS 0.181057f
C2458 vernier_delay_line_0.stop_strong.t1 VSS 0.055955f
C2459 vernier_delay_line_0.stop_strong.n17 VSS 0.413796f
C2460 vernier_delay_line_0.stop_strong.n18 VSS 0.11234f
C2461 vernier_delay_line_0.stop_strong.t10 VSS 0.181057f
C2462 vernier_delay_line_0.stop_strong.t11 VSS 0.055955f
C2463 vernier_delay_line_0.stop_strong.n19 VSS 0.413796f
C2464 vernier_delay_line_0.stop_strong.n20 VSS 0.11234f
C2465 vernier_delay_line_0.stop_strong.t31 VSS 0.181057f
C2466 vernier_delay_line_0.stop_strong.t22 VSS 0.055955f
C2467 vernier_delay_line_0.stop_strong.n21 VSS 0.413796f
C2468 vernier_delay_line_0.stop_strong.n22 VSS 0.11234f
C2469 vernier_delay_line_0.stop_strong.t24 VSS 0.181057f
C2470 vernier_delay_line_0.stop_strong.t25 VSS 0.055955f
C2471 vernier_delay_line_0.stop_strong.n23 VSS 0.413796f
C2472 vernier_delay_line_0.stop_strong.n24 VSS 0.11234f
C2473 vernier_delay_line_0.stop_strong.t13 VSS 0.181057f
C2474 vernier_delay_line_0.stop_strong.t17 VSS 0.055955f
C2475 vernier_delay_line_0.stop_strong.n25 VSS 0.413796f
C2476 vernier_delay_line_0.stop_strong.n26 VSS 0.11234f
C2477 vernier_delay_line_0.stop_strong.t5 VSS 0.181057f
C2478 vernier_delay_line_0.stop_strong.t30 VSS 0.055955f
C2479 vernier_delay_line_0.stop_strong.n27 VSS 0.413796f
C2480 vernier_delay_line_0.stop_strong.n28 VSS 0.11234f
C2481 vernier_delay_line_0.stop_strong.t23 VSS 0.181057f
C2482 vernier_delay_line_0.stop_strong.t29 VSS 0.055955f
C2483 vernier_delay_line_0.stop_strong.n29 VSS 0.413796f
C2484 vernier_delay_line_0.stop_strong.n30 VSS 0.11234f
C2485 vernier_delay_line_0.stop_strong.t19 VSS 0.181057f
C2486 vernier_delay_line_0.stop_strong.t12 VSS 0.055955f
C2487 vernier_delay_line_0.stop_strong.n31 VSS 0.413796f
C2488 vernier_delay_line_0.stop_strong.n32 VSS 0.11234f
C2489 vernier_delay_line_0.stop_strong.t7 VSS 0.181057f
C2490 vernier_delay_line_0.stop_strong.t4 VSS 0.055955f
C2491 vernier_delay_line_0.stop_strong.n33 VSS 0.413796f
C2492 vernier_delay_line_0.stop_strong.n34 VSS 0.110532f
C2493 vernier_delay_line_0.stop_strong.t26 VSS 0.179153f
C2494 vernier_delay_line_0.stop_strong.t27 VSS 0.055955f
C2495 vernier_delay_line_0.stop_strong.n35 VSS 1.27701f
C2496 vernier_delay_line_0.saff_delay_unit_0/saff_2_0.sense_amplifier_0.clk VSS 0.970791f
C2497 vernier_delay_line_0.stop_strong.t64 VSS 0.093756f
C2498 vernier_delay_line_0.stop_strong.t50 VSS 0.093545f
C2499 vernier_delay_line_0.stop_strong.n36 VSS 0.403473f
C2500 vernier_delay_line_0.stop_strong.t42 VSS 0.072027f
C2501 vernier_delay_line_0.stop_strong.t58 VSS 0.072027f
C2502 vernier_delay_line_0.stop_strong.t34 VSS 0.072027f
C2503 vernier_delay_line_0.stop_strong.t39 VSS 0.072027f
C2504 vernier_delay_line_0.stop_strong.t65 VSS 0.079805f
C2505 vernier_delay_line_0.stop_strong.n37 VSS 0.070183f
C2506 vernier_delay_line_0.stop_strong.n38 VSS 0.04137f
C2507 vernier_delay_line_0.stop_strong.n39 VSS 0.04137f
C2508 vernier_delay_line_0.stop_strong.n40 VSS 0.062319f
C2509 vernier_delay_line_0.stop_strong.n41 VSS 0.781253f
C2510 vernier_delay_line_0.stop_strong.n42 VSS 0.697924f
C2511 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2512 vernier_delay_line_0.stop_strong.t74 VSS 0.093756f
C2513 vernier_delay_line_0.stop_strong.t77 VSS 0.093545f
C2514 vernier_delay_line_0.stop_strong.n43 VSS 0.403473f
C2515 vernier_delay_line_0.stop_strong.t57 VSS 0.072027f
C2516 vernier_delay_line_0.stop_strong.t33 VSS 0.072027f
C2517 vernier_delay_line_0.stop_strong.t47 VSS 0.072027f
C2518 vernier_delay_line_0.stop_strong.t70 VSS 0.072027f
C2519 vernier_delay_line_0.stop_strong.t36 VSS 0.079805f
C2520 vernier_delay_line_0.stop_strong.n44 VSS 0.070183f
C2521 vernier_delay_line_0.stop_strong.n45 VSS 0.04137f
C2522 vernier_delay_line_0.stop_strong.n46 VSS 0.04137f
C2523 vernier_delay_line_0.stop_strong.n47 VSS 0.062319f
C2524 vernier_delay_line_0.stop_strong.n48 VSS 0.781253f
C2525 vernier_delay_line_0.stop_strong.n49 VSS 0.697924f
C2526 vernier_delay_line_0.saff_delay_unit_2/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2527 vernier_delay_line_0.stop_strong.t85 VSS 0.093756f
C2528 vernier_delay_line_0.stop_strong.t45 VSS 0.093545f
C2529 vernier_delay_line_0.stop_strong.n50 VSS 0.403473f
C2530 vernier_delay_line_0.stop_strong.t78 VSS 0.072027f
C2531 vernier_delay_line_0.stop_strong.t46 VSS 0.072027f
C2532 vernier_delay_line_0.stop_strong.t69 VSS 0.072027f
C2533 vernier_delay_line_0.stop_strong.t35 VSS 0.072027f
C2534 vernier_delay_line_0.stop_strong.t49 VSS 0.079805f
C2535 vernier_delay_line_0.stop_strong.n51 VSS 0.070183f
C2536 vernier_delay_line_0.stop_strong.n52 VSS 0.04137f
C2537 vernier_delay_line_0.stop_strong.n53 VSS 0.04137f
C2538 vernier_delay_line_0.stop_strong.n54 VSS 0.062319f
C2539 vernier_delay_line_0.stop_strong.n55 VSS 0.781253f
C2540 vernier_delay_line_0.stop_strong.n56 VSS 0.697924f
C2541 vernier_delay_line_0.saff_delay_unit_3/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2542 vernier_delay_line_0.stop_strong.t56 VSS 0.093756f
C2543 vernier_delay_line_0.stop_strong.t60 VSS 0.093545f
C2544 vernier_delay_line_0.stop_strong.n57 VSS 0.403473f
C2545 vernier_delay_line_0.stop_strong.t53 VSS 0.072027f
C2546 vernier_delay_line_0.stop_strong.t61 VSS 0.072027f
C2547 vernier_delay_line_0.stop_strong.t81 VSS 0.072027f
C2548 vernier_delay_line_0.stop_strong.t48 VSS 0.072027f
C2549 vernier_delay_line_0.stop_strong.t87 VSS 0.079805f
C2550 vernier_delay_line_0.stop_strong.n58 VSS 0.070183f
C2551 vernier_delay_line_0.stop_strong.n59 VSS 0.04137f
C2552 vernier_delay_line_0.stop_strong.n60 VSS 0.04137f
C2553 vernier_delay_line_0.stop_strong.n61 VSS 0.062319f
C2554 vernier_delay_line_0.stop_strong.n62 VSS 0.781253f
C2555 vernier_delay_line_0.stop_strong.n63 VSS 0.697924f
C2556 vernier_delay_line_0.saff_delay_unit_4/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2557 vernier_delay_line_0.stop_strong.t71 VSS 0.093756f
C2558 vernier_delay_line_0.stop_strong.t68 VSS 0.093545f
C2559 vernier_delay_line_0.stop_strong.n64 VSS 0.403473f
C2560 vernier_delay_line_0.stop_strong.t52 VSS 0.072027f
C2561 vernier_delay_line_0.stop_strong.t73 VSS 0.072027f
C2562 vernier_delay_line_0.stop_strong.t41 VSS 0.072027f
C2563 vernier_delay_line_0.stop_strong.t82 VSS 0.072027f
C2564 vernier_delay_line_0.stop_strong.t86 VSS 0.079805f
C2565 vernier_delay_line_0.stop_strong.n65 VSS 0.070183f
C2566 vernier_delay_line_0.stop_strong.n66 VSS 0.04137f
C2567 vernier_delay_line_0.stop_strong.n67 VSS 0.04137f
C2568 vernier_delay_line_0.stop_strong.n68 VSS 0.062319f
C2569 vernier_delay_line_0.stop_strong.n69 VSS 0.781253f
C2570 vernier_delay_line_0.stop_strong.n70 VSS 0.697924f
C2571 vernier_delay_line_0.saff_delay_unit_5/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2572 vernier_delay_line_0.stop_strong.t37 VSS 0.093756f
C2573 vernier_delay_line_0.stop_strong.t40 VSS 0.093545f
C2574 vernier_delay_line_0.stop_strong.n71 VSS 0.403473f
C2575 vernier_delay_line_0.stop_strong.t63 VSS 0.072027f
C2576 vernier_delay_line_0.stop_strong.t84 VSS 0.072027f
C2577 vernier_delay_line_0.stop_strong.t66 VSS 0.072027f
C2578 vernier_delay_line_0.stop_strong.t32 VSS 0.072027f
C2579 vernier_delay_line_0.stop_strong.t62 VSS 0.079805f
C2580 vernier_delay_line_0.stop_strong.n72 VSS 0.070183f
C2581 vernier_delay_line_0.stop_strong.n73 VSS 0.04137f
C2582 vernier_delay_line_0.stop_strong.n74 VSS 0.04137f
C2583 vernier_delay_line_0.stop_strong.n75 VSS 0.062319f
C2584 vernier_delay_line_0.stop_strong.n76 VSS 0.781253f
C2585 vernier_delay_line_0.stop_strong.n77 VSS 0.697924f
C2586 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.clk VSS 0.626873f
C2587 vernier_delay_line_0.stop_strong.t51 VSS 0.093756f
C2588 vernier_delay_line_0.stop_strong.t54 VSS 0.093545f
C2589 vernier_delay_line_0.stop_strong.n78 VSS 0.403473f
C2590 vernier_delay_line_0.stop_strong.t83 VSS 0.072027f
C2591 vernier_delay_line_0.stop_strong.t55 VSS 0.072027f
C2592 vernier_delay_line_0.stop_strong.t76 VSS 0.072027f
C2593 vernier_delay_line_0.stop_strong.t44 VSS 0.072027f
C2594 vernier_delay_line_0.stop_strong.t67 VSS 0.079805f
C2595 vernier_delay_line_0.stop_strong.n79 VSS 0.070183f
C2596 vernier_delay_line_0.stop_strong.n80 VSS 0.04137f
C2597 vernier_delay_line_0.stop_strong.n81 VSS 0.04137f
C2598 vernier_delay_line_0.stop_strong.n82 VSS 0.062319f
C2599 vernier_delay_line_0.stop_strong.n83 VSS 0.781253f
C2600 vernier_delay_line_0.stop_strong.n84 VSS 0.697924f
C2601 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.clk VSS 1.31509f
C2602 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C2603 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C2604 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.087567f
C2605 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.039891f
C2606 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C2607 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.201734f
C2608 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C2609 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.095888f
C2610 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.041221f
C2611 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C2612 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.108538f
C2613 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.081767f
C2614 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.090596f
C2615 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C2616 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C2617 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C2618 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C2619 vernier_delay_line_0.saff_delay_unit_1/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C2620 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C2621 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C2622 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.087567f
C2623 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.039891f
C2624 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C2625 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.201734f
C2626 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.201734f
C2627 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.095888f
C2628 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.041221f
C2629 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.116123f
C2630 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.108538f
C2631 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.081767f
C2632 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.090596f
C2633 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.106694f
C2634 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.054262f
C2635 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.054262f
C2636 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.115133f
C2637 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C2638 diff_gen_0.delay_unit_2_6.in_1.t13 VSS 0.086195f
C2639 diff_gen_0.delay_unit_2_6.in_1.t8 VSS 0.027496f
C2640 diff_gen_0.delay_unit_2_6.in_1.n0 VSS 0.060063f
C2641 diff_gen_0.delay_unit_2_6.in_1.t10 VSS 0.086195f
C2642 diff_gen_0.delay_unit_2_6.in_1.t11 VSS 0.027496f
C2643 diff_gen_0.delay_unit_2_6.in_1.n1 VSS 0.060453f
C2644 diff_gen_0.delay_unit_2_6.in_1.n2 VSS 0.019374f
C2645 diff_gen_0.delay_unit_2_6.in_1.t14 VSS 0.086195f
C2646 diff_gen_0.delay_unit_2_6.in_1.t9 VSS 0.027496f
C2647 diff_gen_0.delay_unit_2_6.in_1.n3 VSS 0.060453f
C2648 diff_gen_0.delay_unit_2_6.in_1.t12 VSS 0.086195f
C2649 diff_gen_0.delay_unit_2_6.in_1.t15 VSS 0.027496f
C2650 diff_gen_0.delay_unit_2_6.in_1.n4 VSS 0.060063f
C2651 diff_gen_0.delay_unit_2_6.in_1.n5 VSS 0.019163f
C2652 diff_gen_0.delay_unit_2_6.in_1.n6 VSS 0.505752f
C2653 diff_gen_0.delay_unit_2_6.in_1.t7 VSS 0.068982f
C2654 diff_gen_0.delay_unit_2_6.in_1.t6 VSS 0.2088f
C2655 diff_gen_0.delay_unit_2_6.in_1.n7 VSS 0.529943f
C2656 diff_gen_0.delay_unit_2_6.in_1.n8 VSS 0.27619f
C2657 diff_gen_0.delay_unit_2_6.in_1.t1 VSS 0.018851f
C2658 diff_gen_0.delay_unit_2_6.in_1.t2 VSS 0.018851f
C2659 diff_gen_0.delay_unit_2_6.in_1.n9 VSS 0.044154f
C2660 diff_gen_0.delay_unit_2_6.in_1.t5 VSS 0.056553f
C2661 diff_gen_0.delay_unit_2_6.in_1.t3 VSS 0.056553f
C2662 diff_gen_0.delay_unit_2_6.in_1.n10 VSS 0.115209f
C2663 diff_gen_0.delay_unit_2_6.in_1.n11 VSS 0.479339f
C2664 diff_gen_0.delay_unit_2_6.in_1.t0 VSS 0.069002f
C2665 diff_gen_0.delay_unit_2_6.in_1.t4 VSS 0.2088f
C2666 diff_gen_0.delay_unit_2_6.in_1.n12 VSS 0.509237f
C2667 diff_gen_0.delay_unit_2_6.in_1.n13 VSS 0.26045f
C2668 diff_gen_0.delay_unit_2_5.in_2.n0 VSS 0.400401f
C2669 diff_gen_0.delay_unit_2_5.in_2.t13 VSS 0.066664f
C2670 diff_gen_0.delay_unit_2_5.in_2.t15 VSS 0.021266f
C2671 diff_gen_0.delay_unit_2_5.in_2.n1 VSS 0.046756f
C2672 diff_gen_0.delay_unit_2_5.in_2.t10 VSS 0.066664f
C2673 diff_gen_0.delay_unit_2_5.in_2.t12 VSS 0.021266f
C2674 diff_gen_0.delay_unit_2_5.in_2.n2 VSS 0.046454f
C2675 diff_gen_0.delay_unit_2_5.in_2.n3 VSS 0.014982f
C2676 diff_gen_0.delay_unit_2_5.in_2.t14 VSS 0.066664f
C2677 diff_gen_0.delay_unit_2_5.in_2.t8 VSS 0.021266f
C2678 diff_gen_0.delay_unit_2_5.in_2.n4 VSS 0.046756f
C2679 diff_gen_0.delay_unit_2_5.in_2.t9 VSS 0.066664f
C2680 diff_gen_0.delay_unit_2_5.in_2.t11 VSS 0.021266f
C2681 diff_gen_0.delay_unit_2_5.in_2.n5 VSS 0.046454f
C2682 diff_gen_0.delay_unit_2_5.in_2.n6 VSS 0.014821f
C2683 diff_gen_0.delay_unit_2_5.in_2.n7 VSS 0.22891f
C2684 diff_gen_0.delay_unit_2_5.in_2.t4 VSS 0.165681f
C2685 diff_gen_0.delay_unit_2_5.in_2.t2 VSS 0.051203f
C2686 diff_gen_0.delay_unit_2_5.in_2.n8 VSS 0.452839f
C2687 diff_gen_0.delay_unit_2_5.in_2.t0 VSS 0.043739f
C2688 diff_gen_0.delay_unit_2_5.in_2.t1 VSS 0.043739f
C2689 diff_gen_0.delay_unit_2_5.in_2.n9 VSS 0.093535f
C2690 diff_gen_0.delay_unit_2_5.in_2.t6 VSS 0.01458f
C2691 diff_gen_0.delay_unit_2_5.in_2.t7 VSS 0.01458f
C2692 diff_gen_0.delay_unit_2_5.in_2.n10 VSS 0.031652f
C2693 diff_gen_0.delay_unit_2_5.in_2.n11 VSS 0.376142f
C2694 diff_gen_0.delay_unit_2_5.in_2.t3 VSS 0.165681f
C2695 diff_gen_0.delay_unit_2_5.in_2.t5 VSS 0.051203f
C2696 diff_gen_0.delay_unit_2_5.in_2.n12 VSS 0.398173f
C2697 a_14774_2192.t3 VSS 0.024913f
C2698 a_14774_2192.t8 VSS 0.024913f
C2699 a_14774_2192.n0 VSS 0.060114f
C2700 a_14774_2192.t7 VSS 0.024913f
C2701 a_14774_2192.t6 VSS 0.024913f
C2702 a_14774_2192.n1 VSS 0.060114f
C2703 a_14774_2192.t4 VSS 0.024913f
C2704 a_14774_2192.t9 VSS 0.024913f
C2705 a_14774_2192.n2 VSS 0.060114f
C2706 a_14774_2192.t1 VSS 0.024913f
C2707 a_14774_2192.t0 VSS 0.024913f
C2708 a_14774_2192.n3 VSS 0.057409f
C2709 a_14774_2192.t5 VSS 0.024913f
C2710 a_14774_2192.t2 VSS 0.024913f
C2711 a_14774_2192.n4 VSS 0.060272f
C2712 a_14774_2192.n5 VSS 0.340434f
C2713 a_14774_2192.t12 VSS 0.024913f
C2714 a_14774_2192.t11 VSS 0.024913f
C2715 a_14774_2192.n6 VSS 0.052659f
C2716 a_14774_2192.n7 VSS 0.140942f
C2717 a_14774_2192.n8 VSS 0.22019f
C2718 a_14774_2192.n9 VSS 0.182473f
C2719 a_14774_2192.n10 VSS 0.369186f
C2720 a_14774_2192.t10 VSS 0.097139f
C2721 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t19 VSS 0.059856f
C2722 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t10 VSS 0.019094f
C2723 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n0 VSS 0.041709f
C2724 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t13 VSS 0.059856f
C2725 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t16 VSS 0.019094f
C2726 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n1 VSS 0.04198f
C2727 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n2 VSS 0.013454f
C2728 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t18 VSS 0.059856f
C2729 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t9 VSS 0.019094f
C2730 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n3 VSS 0.04198f
C2731 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t11 VSS 0.059856f
C2732 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t14 VSS 0.019094f
C2733 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n4 VSS 0.041709f
C2734 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n5 VSS 0.013307f
C2735 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n6 VSS 0.351208f
C2736 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t4 VSS 0.047903f
C2737 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t5 VSS 0.144997f
C2738 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n7 VSS 0.368007f
C2739 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t7 VSS 0.013091f
C2740 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t2 VSS 0.013091f
C2741 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n8 VSS 0.030662f
C2742 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t1 VSS 0.039272f
C2743 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t0 VSS 0.039272f
C2744 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n9 VSS 0.080004f
C2745 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n10 VSS 0.332866f
C2746 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t12 VSS 0.061472f
C2747 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t17 VSS 0.061472f
C2748 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n11 VSS 0.069399f
C2749 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t15 VSS 0.061472f
C2750 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t8 VSS 0.061472f
C2751 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n12 VSS 0.069022f
C2752 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n13 VSS 0.63019f
C2753 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t3 VSS 0.045973f
C2754 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n14 VSS 0.158781f
C2755 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.t6 VSS 0.144997f
C2756 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n15 VSS 0.240639f
C2757 vernier_delay_line_0.saff_delay_unit_7/delay_unit_2_0.in_1.n16 VSS 0.180864f
C2758 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C2759 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.087824f
C2760 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.040008f
C2761 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.097717f
C2762 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.200111f
C2763 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.202807f
C2764 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.096169f
C2765 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.041341f
C2766 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.116331f
C2767 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.082007f
C2768 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.090862f
C2769 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.108213f
C2770 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n4 VSS 1.24645f
C2771 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.107599f
C2772 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C2773 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C2774 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.054421f
C2775 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.114315f
C2776 vernier_delay_line_0.saff_delay_unit_7/saff_2_0.sense_amplifier_0.out1.n7 VSS 0.382243f
C2777 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n0 VSS 0.763336f
C2778 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n1 VSS 0.936187f
C2779 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t5 VSS 0.087567f
C2780 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t10 VSS 0.039891f
C2781 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n2 VSS 0.097546f
C2782 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t3 VSS 0.054262f
C2783 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t2 VSS 0.054262f
C2784 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n3 VSS 0.115133f
C2785 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t1 VSS 0.201734f
C2786 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t7 VSS 0.095888f
C2787 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t6 VSS 0.041221f
C2788 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n4 VSS 0.116123f
C2789 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t9 VSS 0.108538f
C2790 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t4 VSS 0.081767f
C2791 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t8 VSS 0.090596f
C2792 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n5 VSS 0.106694f
C2793 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.t0 VSS 0.201734f
C2794 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out2.n6 VSS 0.753756f
C2795 VDD.n0 VSS 0.100844f
C2796 VDD.t223 VSS 0.019607f
C2797 VDD.t406 VSS 0.019607f
C2798 VDD.n1 VSS 0.04155f
C2799 VDD.t219 VSS 0.073915f
C2800 VDD.n2 VSS 0.071633f
C2801 VDD.t29 VSS 0.073915f
C2802 VDD.n3 VSS 0.170163f
C2803 VDD.t87 VSS 0.019607f
C2804 VDD.t503 VSS 0.019607f
C2805 VDD.n4 VSS 0.04155f
C2806 VDD.n5 VSS 0.356059f
C2807 VDD.n6 VSS 0.119907f
C2808 VDD.n7 VSS 0.387327f
C2809 VDD.n8 VSS 0.146538f
C2810 VDD.t86 VSS 0.301845f
C2811 VDD.t502 VSS 0.190393f
C2812 VDD.t495 VSS 0.190393f
C2813 VDD.t28 VSS 0.249891f
C2814 VDD.n9 VSS 0.383723f
C2815 VDD.t405 VSS 0.296651f
C2816 VDD.t222 VSS 0.190393f
C2817 VDD.t197 VSS 0.190393f
C2818 VDD.t218 VSS 0.252054f
C2819 VDD.n10 VSS 0.043203f
C2820 VDD.n11 VSS 0.159021f
C2821 VDD.n12 VSS 0.156858f
C2822 VDD.n13 VSS 0.129206f
C2823 VDD.n14 VSS 0.146538f
C2824 VDD.n15 VSS 0.129206f
C2825 VDD.n16 VSS 0.011609f
C2826 VDD.n17 VSS 0.064542f
C2827 VDD.n18 VSS 0.170393f
C2828 VDD.n19 VSS 0.173658f
C2829 VDD.n20 VSS 0.085001f
C2830 VDD.n21 VSS 0.100989f
C2831 VDD.t363 VSS 0.019607f
C2832 VDD.t439 VSS 0.019607f
C2833 VDD.n22 VSS 0.04155f
C2834 VDD.t83 VSS 0.073915f
C2835 VDD.n23 VSS 0.064542f
C2836 VDD.n24 VSS 0.129206f
C2837 VDD.n25 VSS 0.071633f
C2838 VDD.t361 VSS 0.019607f
C2839 VDD.t367 VSS 0.019607f
C2840 VDD.n26 VSS 0.04155f
C2841 VDD.t435 VSS 0.073915f
C2842 VDD.n27 VSS 0.170393f
C2843 VDD.n28 VSS 0.173658f
C2844 VDD.n29 VSS 0.100989f
C2845 VDD.t329 VSS 0.019607f
C2846 VDD.t59 VSS 0.019607f
C2847 VDD.n30 VSS 0.04155f
C2848 VDD.t128 VSS 0.073915f
C2849 VDD.n31 VSS 0.064542f
C2850 VDD.n32 VSS 0.129206f
C2851 VDD.n33 VSS 0.071633f
C2852 VDD.t392 VSS 0.019607f
C2853 VDD.t390 VSS 0.019607f
C2854 VDD.n34 VSS 0.04155f
C2855 VDD.t384 VSS 0.073915f
C2856 VDD.n35 VSS 0.170393f
C2857 VDD.n36 VSS 0.173658f
C2858 VDD.n37 VSS 0.100989f
C2859 VDD.t420 VSS 0.019607f
C2860 VDD.t422 VSS 0.019607f
C2861 VDD.n38 VSS 0.04155f
C2862 VDD.t25 VSS 0.073915f
C2863 VDD.n39 VSS 0.064542f
C2864 VDD.n40 VSS 0.129206f
C2865 VDD.n41 VSS 0.071633f
C2866 VDD.t426 VSS 0.019607f
C2867 VDD.t428 VSS 0.019607f
C2868 VDD.n42 VSS 0.04155f
C2869 VDD.t155 VSS 0.073915f
C2870 VDD.n43 VSS 0.170393f
C2871 VDD.n44 VSS 0.173658f
C2872 VDD.n45 VSS 0.100989f
C2873 VDD.t1 VSS 0.019607f
C2874 VDD.t140 VSS 0.019607f
C2875 VDD.n46 VSS 0.04155f
C2876 VDD.t470 VSS 0.073915f
C2877 VDD.n47 VSS 0.064542f
C2878 VDD.n48 VSS 0.129206f
C2879 VDD.n49 VSS 0.071633f
C2880 VDD.t5 VSS 0.019607f
C2881 VDD.t142 VSS 0.019607f
C2882 VDD.n50 VSS 0.04155f
C2883 VDD.t388 VSS 0.073915f
C2884 VDD.n51 VSS 0.170393f
C2885 VDD.n52 VSS 0.173658f
C2886 VDD.n53 VSS 0.100989f
C2887 VDD.t445 VSS 0.019607f
C2888 VDD.t138 VSS 0.019607f
C2889 VDD.n54 VSS 0.04155f
C2890 VDD.t287 VSS 0.073915f
C2891 VDD.n55 VSS 0.064542f
C2892 VDD.n56 VSS 0.129206f
C2893 VDD.n57 VSS 0.071633f
C2894 VDD.t459 VSS 0.019607f
C2895 VDD.t275 VSS 0.019607f
C2896 VDD.n58 VSS 0.04155f
C2897 VDD.t194 VSS 0.073915f
C2898 VDD.n59 VSS 0.170393f
C2899 VDD.n60 VSS 0.173658f
C2900 VDD.n61 VSS 0.100989f
C2901 VDD.t343 VSS 0.019607f
C2902 VDD.t398 VSS 0.019607f
C2903 VDD.n62 VSS 0.04155f
C2904 VDD.t157 VSS 0.073915f
C2905 VDD.n63 VSS 0.064542f
C2906 VDD.n64 VSS 0.129206f
C2907 VDD.n65 VSS 0.071633f
C2908 VDD.t226 VSS 0.019607f
C2909 VDD.t136 VSS 0.019607f
C2910 VDD.n66 VSS 0.04155f
C2911 VDD.t271 VSS 0.073915f
C2912 VDD.n67 VSS 0.170393f
C2913 VDD.n68 VSS 0.173658f
C2914 VDD.n69 VSS 0.100989f
C2915 VDD.t297 VSS 0.019607f
C2916 VDD.t261 VSS 0.019607f
C2917 VDD.n70 VSS 0.04155f
C2918 VDD.t190 VSS 0.073915f
C2919 VDD.n71 VSS 0.064542f
C2920 VDD.n72 VSS 0.129206f
C2921 VDD.n73 VSS 0.071633f
C2922 VDD.t291 VSS 0.019607f
C2923 VDD.t349 VSS 0.019607f
C2924 VDD.n74 VSS 0.04155f
C2925 VDD.t234 VSS 0.073915f
C2926 VDD.n75 VSS 0.170393f
C2927 VDD.n76 VSS 0.173658f
C2928 VDD.n77 VSS 0.298764f
C2929 VDD.t447 VSS 0.073581f
C2930 VDD.n78 VSS 0.135752f
C2931 VDD.n79 VSS 0.06005f
C2932 VDD.n80 VSS 0.063491f
C2933 VDD.n81 VSS 0.031372f
C2934 VDD.n82 VSS 0.045083f
C2935 VDD.n83 VSS 0.075491f
C2936 VDD.t91 VSS 0.073581f
C2937 VDD.n84 VSS 0.063491f
C2938 VDD.t267 VSS 0.073581f
C2939 VDD.n85 VSS 0.135752f
C2940 VDD.n86 VSS 0.031372f
C2941 VDD.n87 VSS 0.063491f
C2942 VDD.n88 VSS 0.031372f
C2943 VDD.n89 VSS 0.045083f
C2944 VDD.n90 VSS 0.075491f
C2945 VDD.t305 VSS 0.073581f
C2946 VDD.n91 VSS 0.063491f
C2947 VDD.t85 VSS 0.073581f
C2948 VDD.n92 VSS 0.135752f
C2949 VDD.n93 VSS 0.031372f
C2950 VDD.n94 VSS 0.063491f
C2951 VDD.n95 VSS 0.031372f
C2952 VDD.n96 VSS 0.045083f
C2953 VDD.n97 VSS 0.075491f
C2954 VDD.t167 VSS 0.073581f
C2955 VDD.n98 VSS 0.063491f
C2956 VDD.t333 VSS 0.073581f
C2957 VDD.n99 VSS 0.135752f
C2958 VDD.n100 VSS 0.031372f
C2959 VDD.n101 VSS 0.063491f
C2960 VDD.n102 VSS 0.031372f
C2961 VDD.n103 VSS 0.045083f
C2962 VDD.n104 VSS 0.075491f
C2963 VDD.t488 VSS 0.073581f
C2964 VDD.n105 VSS 0.063491f
C2965 VDD.t109 VSS 0.073581f
C2966 VDD.n106 VSS 0.135752f
C2967 VDD.n107 VSS 0.031372f
C2968 VDD.n108 VSS 0.063491f
C2969 VDD.n109 VSS 0.031372f
C2970 VDD.n110 VSS 0.045083f
C2971 VDD.n111 VSS 0.075491f
C2972 VDD.t7 VSS 0.073581f
C2973 VDD.n112 VSS 0.063491f
C2974 VDD.t169 VSS 0.073581f
C2975 VDD.n113 VSS 0.135752f
C2976 VDD.n114 VSS 0.031372f
C2977 VDD.n115 VSS 0.063491f
C2978 VDD.n116 VSS 0.031372f
C2979 VDD.n117 VSS 0.045083f
C2980 VDD.n118 VSS 0.075491f
C2981 VDD.t89 VSS 0.073581f
C2982 VDD.n119 VSS 0.063491f
C2983 VDD.t265 VSS 0.073581f
C2984 VDD.n120 VSS 0.135752f
C2985 VDD.n121 VSS 0.031372f
C2986 VDD.n122 VSS 0.063491f
C2987 VDD.n123 VSS 0.031372f
C2988 VDD.n124 VSS 0.045083f
C2989 VDD.n125 VSS 0.075491f
C2990 VDD.t43 VSS 0.073581f
C2991 VDD.n126 VSS 0.063491f
C2992 VDD.t107 VSS 0.073581f
C2993 VDD.n127 VSS 0.135752f
C2994 VDD.n128 VSS 0.031372f
C2995 VDD.n129 VSS 0.063491f
C2996 VDD.n130 VSS 0.031372f
C2997 VDD.n131 VSS 0.045083f
C2998 VDD.n132 VSS 0.075491f
C2999 VDD.t303 VSS 0.073581f
C3000 VDD.n133 VSS 0.063491f
C3001 VDD.t203 VSS 0.073581f
C3002 VDD.n134 VSS 0.135752f
C3003 VDD.n135 VSS 0.031372f
C3004 VDD.n136 VSS 0.063491f
C3005 VDD.n137 VSS 0.031372f
C3006 VDD.n138 VSS 0.045083f
C3007 VDD.n139 VSS 0.075491f
C3008 VDD.t199 VSS 0.073581f
C3009 VDD.n140 VSS 0.063491f
C3010 VDD.t205 VSS 0.073581f
C3011 VDD.n141 VSS 0.135752f
C3012 VDD.n142 VSS 0.031372f
C3013 VDD.n143 VSS 0.063491f
C3014 VDD.n144 VSS 0.031372f
C3015 VDD.n145 VSS 0.045083f
C3016 VDD.n146 VSS 0.075491f
C3017 VDD.t201 VSS 0.073581f
C3018 VDD.n147 VSS 0.063491f
C3019 VDD.t53 VSS 0.073581f
C3020 VDD.n148 VSS 0.135752f
C3021 VDD.n149 VSS 0.031372f
C3022 VDD.n150 VSS 0.063491f
C3023 VDD.n151 VSS 0.031372f
C3024 VDD.n152 VSS 0.045083f
C3025 VDD.n153 VSS 0.075491f
C3026 VDD.t14 VSS 0.073581f
C3027 VDD.n154 VSS 0.063491f
C3028 VDD.t163 VSS 0.073581f
C3029 VDD.n155 VSS 0.135752f
C3030 VDD.n156 VSS 0.031372f
C3031 VDD.n157 VSS 0.063491f
C3032 VDD.n158 VSS 0.031372f
C3033 VDD.n159 VSS 0.045083f
C3034 VDD.n160 VSS 0.075491f
C3035 VDD.t241 VSS 0.073581f
C3036 VDD.n161 VSS 0.063491f
C3037 VDD.t124 VSS 0.073581f
C3038 VDD.n162 VSS 0.135752f
C3039 VDD.n163 VSS 0.031372f
C3040 VDD.n164 VSS 0.063491f
C3041 VDD.n165 VSS 0.031372f
C3042 VDD.n166 VSS 0.045083f
C3043 VDD.n167 VSS 0.075491f
C3044 VDD.t285 VSS 0.073581f
C3045 VDD.n168 VSS 0.063491f
C3046 VDD.t408 VSS 0.073581f
C3047 VDD.n169 VSS 0.135752f
C3048 VDD.n170 VSS 0.031372f
C3049 VDD.n171 VSS 0.063491f
C3050 VDD.n172 VSS 0.06005f
C3051 VDD.n173 VSS 0.030675f
C3052 VDD.t446 VSS 0.307371f
C3053 VDD.n174 VSS 0.045083f
C3054 VDD.n175 VSS 0.040323f
C3055 VDD.n176 VSS 0.27973f
C3056 VDD.t90 VSS 0.27973f
C3057 VDD.n177 VSS 0.045083f
C3058 VDD.n178 VSS 0.040323f
C3059 VDD.n179 VSS 0.27973f
C3060 VDD.t266 VSS 0.27973f
C3061 VDD.n180 VSS 0.045083f
C3062 VDD.n181 VSS 0.040323f
C3063 VDD.n182 VSS 0.27973f
C3064 VDD.t304 VSS 0.27973f
C3065 VDD.n183 VSS 0.045083f
C3066 VDD.n184 VSS 0.040323f
C3067 VDD.n185 VSS 0.27973f
C3068 VDD.t84 VSS 0.27973f
C3069 VDD.n186 VSS 0.045083f
C3070 VDD.n187 VSS 0.040323f
C3071 VDD.n188 VSS 0.27973f
C3072 VDD.t166 VSS 0.27973f
C3073 VDD.n189 VSS 0.045083f
C3074 VDD.n190 VSS 0.040323f
C3075 VDD.n191 VSS 0.27973f
C3076 VDD.t332 VSS 0.27973f
C3077 VDD.n192 VSS 0.045083f
C3078 VDD.n193 VSS 0.040323f
C3079 VDD.n194 VSS 0.27973f
C3080 VDD.t487 VSS 0.27973f
C3081 VDD.n195 VSS 0.045083f
C3082 VDD.n196 VSS 0.040323f
C3083 VDD.n197 VSS 0.27973f
C3084 VDD.t108 VSS 0.27973f
C3085 VDD.n198 VSS 0.045083f
C3086 VDD.n199 VSS 0.040323f
C3087 VDD.n200 VSS 0.27973f
C3088 VDD.t6 VSS 0.27973f
C3089 VDD.n201 VSS 0.045083f
C3090 VDD.n202 VSS 0.040323f
C3091 VDD.n203 VSS 0.27973f
C3092 VDD.t168 VSS 0.27973f
C3093 VDD.n204 VSS 0.045083f
C3094 VDD.n205 VSS 0.040323f
C3095 VDD.n206 VSS 0.27973f
C3096 VDD.t88 VSS 0.27973f
C3097 VDD.n207 VSS 0.045083f
C3098 VDD.n208 VSS 0.040323f
C3099 VDD.n209 VSS 0.27973f
C3100 VDD.t264 VSS 0.27973f
C3101 VDD.n210 VSS 0.045083f
C3102 VDD.n211 VSS 0.040323f
C3103 VDD.n212 VSS 0.27973f
C3104 VDD.t42 VSS 0.27973f
C3105 VDD.n213 VSS 0.045083f
C3106 VDD.n214 VSS 0.040323f
C3107 VDD.n215 VSS 0.27973f
C3108 VDD.t106 VSS 0.27973f
C3109 VDD.n216 VSS 0.045083f
C3110 VDD.n217 VSS 0.040323f
C3111 VDD.n218 VSS 0.27973f
C3112 VDD.t302 VSS 0.27973f
C3113 VDD.n219 VSS 0.045083f
C3114 VDD.n220 VSS 0.040323f
C3115 VDD.n221 VSS 0.27973f
C3116 VDD.t202 VSS 0.27973f
C3117 VDD.n222 VSS 0.045083f
C3118 VDD.n223 VSS 0.040323f
C3119 VDD.n224 VSS 0.27973f
C3120 VDD.t198 VSS 0.27973f
C3121 VDD.n225 VSS 0.045083f
C3122 VDD.n226 VSS 0.040323f
C3123 VDD.n227 VSS 0.27973f
C3124 VDD.t204 VSS 0.27973f
C3125 VDD.n228 VSS 0.045083f
C3126 VDD.n229 VSS 0.040323f
C3127 VDD.n230 VSS 0.27973f
C3128 VDD.t200 VSS 0.27973f
C3129 VDD.n231 VSS 0.045083f
C3130 VDD.n232 VSS 0.040323f
C3131 VDD.n233 VSS 0.27973f
C3132 VDD.t52 VSS 0.27973f
C3133 VDD.n234 VSS 0.045083f
C3134 VDD.n235 VSS 0.040323f
C3135 VDD.n236 VSS 0.27973f
C3136 VDD.t13 VSS 0.27973f
C3137 VDD.n237 VSS 0.045083f
C3138 VDD.n238 VSS 0.040323f
C3139 VDD.n239 VSS 0.27973f
C3140 VDD.t162 VSS 0.27973f
C3141 VDD.n240 VSS 0.045083f
C3142 VDD.n241 VSS 0.040323f
C3143 VDD.n242 VSS 0.27973f
C3144 VDD.t240 VSS 0.27973f
C3145 VDD.n243 VSS 0.045083f
C3146 VDD.n244 VSS 0.040323f
C3147 VDD.n245 VSS 0.27973f
C3148 VDD.t123 VSS 0.27973f
C3149 VDD.n246 VSS 0.045083f
C3150 VDD.n247 VSS 0.040323f
C3151 VDD.n248 VSS 0.27973f
C3152 VDD.t284 VSS 0.27973f
C3153 VDD.n249 VSS 0.045083f
C3154 VDD.n250 VSS 0.040323f
C3155 VDD.n251 VSS 0.27973f
C3156 VDD.t407 VSS 0.27973f
C3157 VDD.n252 VSS 0.045083f
C3158 VDD.n253 VSS 0.040323f
C3159 VDD.n254 VSS 0.27973f
C3160 VDD.t160 VSS 0.307371f
C3161 VDD.n255 VSS 0.030675f
C3162 VDD.n256 VSS 0.298764f
C3163 VDD.n257 VSS 0.075491f
C3164 VDD.t161 VSS 0.073581f
C3165 VDD.n258 VSS 0.065647f
C3166 VDD.n259 VSS 0.135752f
C3167 VDD.n260 VSS 0.020446f
C3168 VDD.n261 VSS 0.06005f
C3169 VDD.n262 VSS 0.045083f
C3170 VDD.n263 VSS 0.031372f
C3171 VDD.n264 VSS 0.020446f
C3172 VDD.n265 VSS 0.075491f
C3173 VDD.n266 VSS 0.135752f
C3174 VDD.n267 VSS 0.020446f
C3175 VDD.n268 VSS 0.031372f
C3176 VDD.n269 VSS 0.045083f
C3177 VDD.n270 VSS 0.031372f
C3178 VDD.n271 VSS 0.020446f
C3179 VDD.n272 VSS 0.075491f
C3180 VDD.n273 VSS 0.135752f
C3181 VDD.n274 VSS 0.020446f
C3182 VDD.n275 VSS 0.031372f
C3183 VDD.n276 VSS 0.045083f
C3184 VDD.n277 VSS 0.031372f
C3185 VDD.n278 VSS 0.020446f
C3186 VDD.n279 VSS 0.075491f
C3187 VDD.n280 VSS 0.135752f
C3188 VDD.n281 VSS 0.020446f
C3189 VDD.n282 VSS 0.031372f
C3190 VDD.n283 VSS 0.045083f
C3191 VDD.n284 VSS 0.031372f
C3192 VDD.n285 VSS 0.020446f
C3193 VDD.n286 VSS 0.075491f
C3194 VDD.n287 VSS 0.135752f
C3195 VDD.n288 VSS 0.020446f
C3196 VDD.n289 VSS 0.031372f
C3197 VDD.n290 VSS 0.045083f
C3198 VDD.n291 VSS 0.031372f
C3199 VDD.n292 VSS 0.020446f
C3200 VDD.n293 VSS 0.075491f
C3201 VDD.n294 VSS 0.135752f
C3202 VDD.n295 VSS 0.020446f
C3203 VDD.n296 VSS 0.031372f
C3204 VDD.n297 VSS 0.045083f
C3205 VDD.n298 VSS 0.031372f
C3206 VDD.n299 VSS 0.020446f
C3207 VDD.n300 VSS 0.075491f
C3208 VDD.n301 VSS 0.135752f
C3209 VDD.n302 VSS 0.020446f
C3210 VDD.n303 VSS 0.031372f
C3211 VDD.n304 VSS 0.045083f
C3212 VDD.n305 VSS 0.031372f
C3213 VDD.n306 VSS 0.020446f
C3214 VDD.n307 VSS 0.075491f
C3215 VDD.n308 VSS 0.135752f
C3216 VDD.n309 VSS 0.020446f
C3217 VDD.n310 VSS 0.031372f
C3218 VDD.n311 VSS 0.045083f
C3219 VDD.n312 VSS 0.031372f
C3220 VDD.n313 VSS 0.020446f
C3221 VDD.n314 VSS 0.075491f
C3222 VDD.n315 VSS 0.135752f
C3223 VDD.n316 VSS 0.020446f
C3224 VDD.n317 VSS 0.031372f
C3225 VDD.n318 VSS 0.045083f
C3226 VDD.n319 VSS 0.031372f
C3227 VDD.n320 VSS 0.020446f
C3228 VDD.n321 VSS 0.075491f
C3229 VDD.n322 VSS 0.135752f
C3230 VDD.n323 VSS 0.020446f
C3231 VDD.n324 VSS 0.031372f
C3232 VDD.n325 VSS 0.045083f
C3233 VDD.n326 VSS 0.031372f
C3234 VDD.n327 VSS 0.020446f
C3235 VDD.n328 VSS 0.075491f
C3236 VDD.n329 VSS 0.135752f
C3237 VDD.n330 VSS 0.020446f
C3238 VDD.n331 VSS 0.031372f
C3239 VDD.n332 VSS 0.045083f
C3240 VDD.n333 VSS 0.031372f
C3241 VDD.n334 VSS 0.020446f
C3242 VDD.n335 VSS 0.075491f
C3243 VDD.n336 VSS 0.135752f
C3244 VDD.n337 VSS 0.020446f
C3245 VDD.n338 VSS 0.031372f
C3246 VDD.n339 VSS 0.045083f
C3247 VDD.n340 VSS 0.031372f
C3248 VDD.n341 VSS 0.020446f
C3249 VDD.n342 VSS 0.075491f
C3250 VDD.n343 VSS 0.135752f
C3251 VDD.n344 VSS 0.020446f
C3252 VDD.n345 VSS 0.031372f
C3253 VDD.n346 VSS 0.045083f
C3254 VDD.n347 VSS 0.031372f
C3255 VDD.n348 VSS 0.020446f
C3256 VDD.n349 VSS 0.075491f
C3257 VDD.n350 VSS 0.135752f
C3258 VDD.n351 VSS 0.020446f
C3259 VDD.n352 VSS 0.031372f
C3260 VDD.n353 VSS 0.045083f
C3261 VDD.n354 VSS 0.06005f
C3262 VDD.n355 VSS 0.020446f
C3263 VDD.n356 VSS 0.143318f
C3264 VDD.n357 VSS 0.100125f
C3265 VDD.t179 VSS 0.07349f
C3266 VDD.t209 VSS 0.07349f
C3267 VDD.t132 VSS 0.07349f
C3268 VDD.t196 VSS 0.074215f
C3269 VDD.n358 VSS 0.27349f
C3270 VDD.n359 VSS 0.145038f
C3271 VDD.n360 VSS 0.135604f
C3272 VDD.n361 VSS 0.100125f
C3273 VDD.t27 VSS 0.07349f
C3274 VDD.t396 VSS 0.07349f
C3275 VDD.t151 VSS 0.07349f
C3276 VDD.t35 VSS 0.074215f
C3277 VDD.n362 VSS 0.27349f
C3278 VDD.n363 VSS 0.145038f
C3279 VDD.n364 VSS 0.135604f
C3280 VDD.n365 VSS 0.100125f
C3281 VDD.t215 VSS 0.07349f
C3282 VDD.t484 VSS 0.07349f
C3283 VDD.t228 VSS 0.07349f
C3284 VDD.t453 VSS 0.074215f
C3285 VDD.n366 VSS 0.27349f
C3286 VDD.n367 VSS 0.145038f
C3287 VDD.n368 VSS 0.135604f
C3288 VDD.n369 VSS 0.100125f
C3289 VDD.t232 VSS 0.07349f
C3290 VDD.t144 VSS 0.07349f
C3291 VDD.t3 VSS 0.07349f
C3292 VDD.t75 VSS 0.074215f
C3293 VDD.n370 VSS 0.27349f
C3294 VDD.n371 VSS 0.145038f
C3295 VDD.n372 VSS 0.135604f
C3296 VDD.n373 VSS 0.100125f
C3297 VDD.t159 VSS 0.07349f
C3298 VDD.t430 VSS 0.07349f
C3299 VDD.t416 VSS 0.07349f
C3300 VDD.t49 VSS 0.074215f
C3301 VDD.n374 VSS 0.27349f
C3302 VDD.n375 VSS 0.145038f
C3303 VDD.n376 VSS 0.135604f
C3304 VDD.n377 VSS 0.100125f
C3305 VDD.t313 VSS 0.07349f
C3306 VDD.t455 VSS 0.07349f
C3307 VDD.t351 VSS 0.07349f
C3308 VDD.t165 VSS 0.074215f
C3309 VDD.n378 VSS 0.27349f
C3310 VDD.n379 VSS 0.145038f
C3311 VDD.n380 VSS 0.135604f
C3312 VDD.n381 VSS 0.100125f
C3313 VDD.t250 VSS 0.07349f
C3314 VDD.t230 VSS 0.07349f
C3315 VDD.t365 VSS 0.07349f
C3316 VDD.t493 VSS 0.074215f
C3317 VDD.n382 VSS 0.27349f
C3318 VDD.n383 VSS 0.145038f
C3319 VDD.n384 VSS 0.135604f
C3320 VDD.n385 VSS 0.100125f
C3321 VDD.t37 VSS 0.07349f
C3322 VDD.t39 VSS 0.07349f
C3323 VDD.t221 VSS 0.07349f
C3324 VDD.t341 VSS 0.074215f
C3325 VDD.n386 VSS 0.27349f
C3326 VDD.n387 VSS 0.145038f
C3327 VDD.n388 VSS 0.135604f
C3328 VDD.n389 VSS 0.458542f
C3329 VDD.n390 VSS 0.412956f
C3330 VDD.t340 VSS 0.318783f
C3331 VDD.t220 VSS 0.352497f
C3332 VDD.n391 VSS 0.263773f
C3333 VDD.n392 VSS 0.33642f
C3334 VDD.t36 VSS 0.314787f
C3335 VDD.t38 VSS 0.369283f
C3336 VDD.n393 VSS 0.722816f
C3337 VDD.n394 VSS 0.069053f
C3338 VDD.n395 VSS 0.694868f
C3339 VDD.n396 VSS 0.384751f
C3340 VDD.n397 VSS 0.157642f
C3341 VDD.n398 VSS 0.458542f
C3342 VDD.n399 VSS 0.412956f
C3343 VDD.t492 VSS 0.318783f
C3344 VDD.t364 VSS 0.352497f
C3345 VDD.n400 VSS 0.263773f
C3346 VDD.n401 VSS 0.33642f
C3347 VDD.t249 VSS 0.314787f
C3348 VDD.t229 VSS 0.369283f
C3349 VDD.n402 VSS 0.722816f
C3350 VDD.n403 VSS 0.069053f
C3351 VDD.n404 VSS 0.455918f
C3352 VDD.n405 VSS 0.299646f
C3353 VDD.n406 VSS 0.089574f
C3354 VDD.n407 VSS 0.157642f
C3355 VDD.n408 VSS 0.458542f
C3356 VDD.n409 VSS 0.412956f
C3357 VDD.t164 VSS 0.318783f
C3358 VDD.t350 VSS 0.352497f
C3359 VDD.n410 VSS 0.263773f
C3360 VDD.n411 VSS 0.33642f
C3361 VDD.t312 VSS 0.314787f
C3362 VDD.t454 VSS 0.369283f
C3363 VDD.n412 VSS 0.722816f
C3364 VDD.n413 VSS 0.069053f
C3365 VDD.n414 VSS 0.455918f
C3366 VDD.n415 VSS 0.299646f
C3367 VDD.n416 VSS 0.089574f
C3368 VDD.n417 VSS 0.157642f
C3369 VDD.n418 VSS 0.458542f
C3370 VDD.n419 VSS 0.412956f
C3371 VDD.t48 VSS 0.318783f
C3372 VDD.t415 VSS 0.352497f
C3373 VDD.n420 VSS 0.263773f
C3374 VDD.n421 VSS 0.33642f
C3375 VDD.t158 VSS 0.314787f
C3376 VDD.t429 VSS 0.369283f
C3377 VDD.n422 VSS 0.722816f
C3378 VDD.n423 VSS 0.069053f
C3379 VDD.n424 VSS 0.455918f
C3380 VDD.n425 VSS 0.299646f
C3381 VDD.n426 VSS 0.089574f
C3382 VDD.n427 VSS 0.157642f
C3383 VDD.n428 VSS 0.458542f
C3384 VDD.n429 VSS 0.412956f
C3385 VDD.t74 VSS 0.318783f
C3386 VDD.t2 VSS 0.352497f
C3387 VDD.n430 VSS 0.263773f
C3388 VDD.n431 VSS 0.33642f
C3389 VDD.t231 VSS 0.314787f
C3390 VDD.t143 VSS 0.369283f
C3391 VDD.n432 VSS 0.722816f
C3392 VDD.n433 VSS 0.069053f
C3393 VDD.n434 VSS 0.455918f
C3394 VDD.n435 VSS 0.299646f
C3395 VDD.n436 VSS 0.089574f
C3396 VDD.n437 VSS 0.157642f
C3397 VDD.n438 VSS 0.458542f
C3398 VDD.n439 VSS 0.412956f
C3399 VDD.t452 VSS 0.318783f
C3400 VDD.t227 VSS 0.352497f
C3401 VDD.n440 VSS 0.263773f
C3402 VDD.n441 VSS 0.33642f
C3403 VDD.t214 VSS 0.314787f
C3404 VDD.t483 VSS 0.369283f
C3405 VDD.n442 VSS 0.722816f
C3406 VDD.n443 VSS 0.069053f
C3407 VDD.n444 VSS 0.455918f
C3408 VDD.n445 VSS 0.299646f
C3409 VDD.n446 VSS 0.089574f
C3410 VDD.n447 VSS 0.157642f
C3411 VDD.n448 VSS 0.458542f
C3412 VDD.n449 VSS 0.412956f
C3413 VDD.t34 VSS 0.318783f
C3414 VDD.t150 VSS 0.352497f
C3415 VDD.n450 VSS 0.263773f
C3416 VDD.n451 VSS 0.33642f
C3417 VDD.t26 VSS 0.314787f
C3418 VDD.t395 VSS 0.369283f
C3419 VDD.n452 VSS 0.722816f
C3420 VDD.n453 VSS 0.069053f
C3421 VDD.n454 VSS 0.455918f
C3422 VDD.n455 VSS 0.299646f
C3423 VDD.n456 VSS 0.089574f
C3424 VDD.n457 VSS 0.157642f
C3425 VDD.n458 VSS 0.458542f
C3426 VDD.n459 VSS 0.412956f
C3427 VDD.t195 VSS 0.318783f
C3428 VDD.t131 VSS 0.352497f
C3429 VDD.n460 VSS 0.263773f
C3430 VDD.n461 VSS 0.33642f
C3431 VDD.t178 VSS 0.314787f
C3432 VDD.t208 VSS 0.369283f
C3433 VDD.n462 VSS 0.722816f
C3434 VDD.n463 VSS 0.069053f
C3435 VDD.n464 VSS 0.455918f
C3436 VDD.n465 VSS 0.299646f
C3437 VDD.n466 VSS 0.089574f
C3438 VDD.n467 VSS 0.157642f
C3439 VDD.n468 VSS 0.114961f
C3440 VDD.t146 VSS 0.019607f
C3441 VDD.t404 VSS 0.019607f
C3442 VDD.n469 VSS 0.041911f
C3443 VDD.t321 VSS 0.019607f
C3444 VDD.t357 VSS 0.019607f
C3445 VDD.n470 VSS 0.041911f
C3446 VDD.t418 VSS 0.019607f
C3447 VDD.t345 VSS 0.019607f
C3448 VDD.n471 VSS 0.041911f
C3449 VDD.n472 VSS 0.168684f
C3450 VDD.n473 VSS 0.138239f
C3451 VDD.n474 VSS 0.11402f
C3452 VDD.t424 VSS 0.019607f
C3453 VDD.t263 VSS 0.019607f
C3454 VDD.n475 VSS 0.041911f
C3455 VDD.n476 VSS 0.169009f
C3456 VDD.n477 VSS 0.090794f
C3457 VDD.t356 VSS 0.268957f
C3458 VDD.t320 VSS 0.202292f
C3459 VDD.t403 VSS 0.202292f
C3460 VDD.t145 VSS 0.300011f
C3461 VDD.n478 VSS 0.335724f
C3462 VDD.n479 VSS 0.132598f
C3463 VDD.n480 VSS 0.100553f
C3464 VDD.n481 VSS 0.172408f
C3465 VDD.n482 VSS 0.167811f
C3466 VDD.t417 VSS 0.264359f
C3467 VDD.t344 VSS 0.202292f
C3468 VDD.t423 VSS 0.202292f
C3469 VDD.t262 VSS 0.267808f
C3470 VDD.t334 VSS 0.267808f
C3471 VDD.n483 VSS 0.132598f
C3472 VDD.n484 VSS 0.138239f
C3473 VDD.t335 VSS 0.019607f
C3474 VDD.t472 VSS 0.019607f
C3475 VDD.n485 VSS 0.041911f
C3476 VDD.t207 VSS 0.019607f
C3477 VDD.t307 VSS 0.019607f
C3478 VDD.n486 VSS 0.041911f
C3479 VDD.t323 VSS 0.019607f
C3480 VDD.t148 VSS 0.019607f
C3481 VDD.n487 VSS 0.041911f
C3482 VDD.n488 VSS 0.168684f
C3483 VDD.n489 VSS 0.11402f
C3484 VDD.t402 VSS 0.019607f
C3485 VDD.t134 VSS 0.019607f
C3486 VDD.n490 VSS 0.041911f
C3487 VDD.n491 VSS 0.169009f
C3488 VDD.n492 VSS 0.090794f
C3489 VDD.t471 VSS 0.202292f
C3490 VDD.t206 VSS 0.202292f
C3491 VDD.t306 VSS 0.268957f
C3492 VDD.n493 VSS 0.100553f
C3493 VDD.n494 VSS 0.172408f
C3494 VDD.n495 VSS 0.167811f
C3495 VDD.t322 VSS 0.264359f
C3496 VDD.t147 VSS 0.202292f
C3497 VDD.t401 VSS 0.202292f
C3498 VDD.t133 VSS 0.267808f
C3499 VDD.t237 VSS 0.267808f
C3500 VDD.n496 VSS 0.132598f
C3501 VDD.n497 VSS 0.138239f
C3502 VDD.t238 VSS 0.019607f
C3503 VDD.t51 VSS 0.019607f
C3504 VDD.n498 VSS 0.041911f
C3505 VDD.t175 VSS 0.019607f
C3506 VDD.t177 VSS 0.019607f
C3507 VDD.n499 VSS 0.041911f
C3508 VDD.t301 VSS 0.019607f
C3509 VDD.t243 VSS 0.019607f
C3510 VDD.n500 VSS 0.041911f
C3511 VDD.n501 VSS 0.168684f
C3512 VDD.n502 VSS 0.11402f
C3513 VDD.t103 VSS 0.019607f
C3514 VDD.t466 VSS 0.019607f
C3515 VDD.n503 VSS 0.041911f
C3516 VDD.n504 VSS 0.169009f
C3517 VDD.n505 VSS 0.090794f
C3518 VDD.t50 VSS 0.202292f
C3519 VDD.t174 VSS 0.202292f
C3520 VDD.t176 VSS 0.268957f
C3521 VDD.n506 VSS 0.100553f
C3522 VDD.n507 VSS 0.172408f
C3523 VDD.n508 VSS 0.167811f
C3524 VDD.t300 VSS 0.264359f
C3525 VDD.t242 VSS 0.202292f
C3526 VDD.t102 VSS 0.202292f
C3527 VDD.t465 VSS 0.267808f
C3528 VDD.t212 VSS 0.267808f
C3529 VDD.n509 VSS 0.132598f
C3530 VDD.n510 VSS 0.138239f
C3531 VDD.t213 VSS 0.019607f
C3532 VDD.t67 VSS 0.019607f
C3533 VDD.n511 VSS 0.041911f
C3534 VDD.t315 VSS 0.019607f
C3535 VDD.t101 VSS 0.019607f
C3536 VDD.n512 VSS 0.041911f
C3537 VDD.t116 VSS 0.019607f
C3538 VDD.t45 VSS 0.019607f
C3539 VDD.n513 VSS 0.041911f
C3540 VDD.n514 VSS 0.168684f
C3541 VDD.n515 VSS 0.11402f
C3542 VDD.t353 VSS 0.019607f
C3543 VDD.t461 VSS 0.019607f
C3544 VDD.n516 VSS 0.041911f
C3545 VDD.n517 VSS 0.169009f
C3546 VDD.n518 VSS 0.090794f
C3547 VDD.t66 VSS 0.202292f
C3548 VDD.t314 VSS 0.202292f
C3549 VDD.t100 VSS 0.268957f
C3550 VDD.n519 VSS 0.100553f
C3551 VDD.n520 VSS 0.172408f
C3552 VDD.n521 VSS 0.167811f
C3553 VDD.t115 VSS 0.264359f
C3554 VDD.t44 VSS 0.202292f
C3555 VDD.t352 VSS 0.202292f
C3556 VDD.t460 VSS 0.267808f
C3557 VDD.t318 VSS 0.267808f
C3558 VDD.n522 VSS 0.132598f
C3559 VDD.n523 VSS 0.138239f
C3560 VDD.t319 VSS 0.019607f
C3561 VDD.t114 VSS 0.019607f
C3562 VDD.n524 VSS 0.041911f
C3563 VDD.t457 VSS 0.019607f
C3564 VDD.t188 VSS 0.019607f
C3565 VDD.n525 VSS 0.041911f
C3566 VDD.t478 VSS 0.019607f
C3567 VDD.t317 VSS 0.019607f
C3568 VDD.n526 VSS 0.041911f
C3569 VDD.n527 VSS 0.168684f
C3570 VDD.n528 VSS 0.11402f
C3571 VDD.t273 VSS 0.019607f
C3572 VDD.t245 VSS 0.019607f
C3573 VDD.n529 VSS 0.041911f
C3574 VDD.n530 VSS 0.169009f
C3575 VDD.n531 VSS 0.090794f
C3576 VDD.t113 VSS 0.202292f
C3577 VDD.t456 VSS 0.202292f
C3578 VDD.t187 VSS 0.268957f
C3579 VDD.n532 VSS 0.100553f
C3580 VDD.n533 VSS 0.172408f
C3581 VDD.n534 VSS 0.167811f
C3582 VDD.t477 VSS 0.264359f
C3583 VDD.t316 VSS 0.202292f
C3584 VDD.t272 VSS 0.202292f
C3585 VDD.t244 VSS 0.267808f
C3586 VDD.t431 VSS 0.267808f
C3587 VDD.n535 VSS 0.132598f
C3588 VDD.n536 VSS 0.138239f
C3589 VDD.t432 VSS 0.019607f
C3590 VDD.t374 VSS 0.019607f
C3591 VDD.n537 VSS 0.041911f
C3592 VDD.t61 VSS 0.019607f
C3593 VDD.t376 VSS 0.019607f
C3594 VDD.n538 VSS 0.041911f
C3595 VDD.t81 VSS 0.019607f
C3596 VDD.t171 VSS 0.019607f
C3597 VDD.n539 VSS 0.041911f
C3598 VDD.n540 VSS 0.168684f
C3599 VDD.n541 VSS 0.11402f
C3600 VDD.t153 VSS 0.019607f
C3601 VDD.t120 VSS 0.019607f
C3602 VDD.n542 VSS 0.041911f
C3603 VDD.n543 VSS 0.169009f
C3604 VDD.n544 VSS 0.090794f
C3605 VDD.t373 VSS 0.202292f
C3606 VDD.t60 VSS 0.202292f
C3607 VDD.t375 VSS 0.268957f
C3608 VDD.n545 VSS 0.100553f
C3609 VDD.n546 VSS 0.172408f
C3610 VDD.n547 VSS 0.167811f
C3611 VDD.t80 VSS 0.264359f
C3612 VDD.t170 VSS 0.202292f
C3613 VDD.t152 VSS 0.202292f
C3614 VDD.t119 VSS 0.267808f
C3615 VDD.t32 VSS 0.267808f
C3616 VDD.n548 VSS 0.132598f
C3617 VDD.n549 VSS 0.138239f
C3618 VDD.t33 VSS 0.019607f
C3619 VDD.t441 VSS 0.019607f
C3620 VDD.n550 VSS 0.041911f
C3621 VDD.t247 VSS 0.019607f
C3622 VDD.t31 VSS 0.019607f
C3623 VDD.n551 VSS 0.041911f
C3624 VDD.t105 VSS 0.019607f
C3625 VDD.t41 VSS 0.019607f
C3626 VDD.n552 VSS 0.041911f
C3627 VDD.n553 VSS 0.168684f
C3628 VDD.n554 VSS 0.11402f
C3629 VDD.t486 VSS 0.019607f
C3630 VDD.t468 VSS 0.019607f
C3631 VDD.n555 VSS 0.041911f
C3632 VDD.n556 VSS 0.169009f
C3633 VDD.n557 VSS 0.298764f
C3634 VDD.t476 VSS 0.073581f
C3635 VDD.n558 VSS 0.135752f
C3636 VDD.n559 VSS 0.06005f
C3637 VDD.n560 VSS 0.063491f
C3638 VDD.n561 VSS 0.031372f
C3639 VDD.n562 VSS 0.045083f
C3640 VDD.n563 VSS 0.075491f
C3641 VDD.t277 VSS 0.073581f
C3642 VDD.n564 VSS 0.063491f
C3643 VDD.t69 VSS 0.073581f
C3644 VDD.n565 VSS 0.135752f
C3645 VDD.n566 VSS 0.031372f
C3646 VDD.n567 VSS 0.063491f
C3647 VDD.n568 VSS 0.031372f
C3648 VDD.n569 VSS 0.045083f
C3649 VDD.n570 VSS 0.075491f
C3650 VDD.t19 VSS 0.073581f
C3651 VDD.n571 VSS 0.063491f
C3652 VDD.t21 VSS 0.073581f
C3653 VDD.n572 VSS 0.135752f
C3654 VDD.n573 VSS 0.031372f
C3655 VDD.n574 VSS 0.063491f
C3656 VDD.n575 VSS 0.031372f
C3657 VDD.n576 VSS 0.045083f
C3658 VDD.n577 VSS 0.075491f
C3659 VDD.t23 VSS 0.073581f
C3660 VDD.n578 VSS 0.063491f
C3661 VDD.t17 VSS 0.073581f
C3662 VDD.n579 VSS 0.135752f
C3663 VDD.n580 VSS 0.031372f
C3664 VDD.n581 VSS 0.063491f
C3665 VDD.n582 VSS 0.06005f
C3666 VDD.n583 VSS 0.030675f
C3667 VDD.t475 VSS 0.307371f
C3668 VDD.n584 VSS 0.045083f
C3669 VDD.n585 VSS 0.040323f
C3670 VDD.n586 VSS 0.27973f
C3671 VDD.t276 VSS 0.27973f
C3672 VDD.n587 VSS 0.045083f
C3673 VDD.n588 VSS 0.040323f
C3674 VDD.n589 VSS 0.27973f
C3675 VDD.t68 VSS 0.27973f
C3676 VDD.n590 VSS 0.045083f
C3677 VDD.n591 VSS 0.040323f
C3678 VDD.n592 VSS 0.27973f
C3679 VDD.t18 VSS 0.27973f
C3680 VDD.n593 VSS 0.045083f
C3681 VDD.n594 VSS 0.040323f
C3682 VDD.n595 VSS 0.27973f
C3683 VDD.t20 VSS 0.27973f
C3684 VDD.n596 VSS 0.045083f
C3685 VDD.n597 VSS 0.040323f
C3686 VDD.n598 VSS 0.27973f
C3687 VDD.t22 VSS 0.27973f
C3688 VDD.n599 VSS 0.045083f
C3689 VDD.n600 VSS 0.040323f
C3690 VDD.n601 VSS 0.27973f
C3691 VDD.t16 VSS 0.27973f
C3692 VDD.n602 VSS 0.045083f
C3693 VDD.n603 VSS 0.040323f
C3694 VDD.n604 VSS 0.27973f
C3695 VDD.t191 VSS 0.307371f
C3696 VDD.n605 VSS 0.030675f
C3697 VDD.n606 VSS 0.298764f
C3698 VDD.n607 VSS 0.075491f
C3699 VDD.t192 VSS 0.073581f
C3700 VDD.n608 VSS 0.065647f
C3701 VDD.n609 VSS 0.135752f
C3702 VDD.n610 VSS 0.020446f
C3703 VDD.n611 VSS 0.06005f
C3704 VDD.n612 VSS 0.045083f
C3705 VDD.n613 VSS 0.031372f
C3706 VDD.n614 VSS 0.020446f
C3707 VDD.n615 VSS 0.075491f
C3708 VDD.n616 VSS 0.135752f
C3709 VDD.n617 VSS 0.020446f
C3710 VDD.n618 VSS 0.031372f
C3711 VDD.n619 VSS 0.045083f
C3712 VDD.n620 VSS 0.031372f
C3713 VDD.n621 VSS 0.020446f
C3714 VDD.n622 VSS 0.075491f
C3715 VDD.n623 VSS 0.135752f
C3716 VDD.n624 VSS 0.020446f
C3717 VDD.n625 VSS 0.031372f
C3718 VDD.n626 VSS 0.045083f
C3719 VDD.n627 VSS 0.031372f
C3720 VDD.n628 VSS 0.020446f
C3721 VDD.n629 VSS 0.075491f
C3722 VDD.n630 VSS 0.135752f
C3723 VDD.n631 VSS 0.020446f
C3724 VDD.n632 VSS 0.031372f
C3725 VDD.n633 VSS 0.045083f
C3726 VDD.n634 VSS 0.06005f
C3727 VDD.n635 VSS 0.020446f
C3728 VDD.n636 VSS 0.100913f
C3729 VDD.n637 VSS 0.084953f
C3730 VDD.t440 VSS 0.202292f
C3731 VDD.t246 VSS 0.202292f
C3732 VDD.t30 VSS 0.268957f
C3733 VDD.n638 VSS 0.100553f
C3734 VDD.n639 VSS 0.172408f
C3735 VDD.n640 VSS 0.167811f
C3736 VDD.t104 VSS 0.264359f
C3737 VDD.t40 VSS 0.202292f
C3738 VDD.t485 VSS 0.202292f
C3739 VDD.t467 VSS 0.267808f
C3740 VDD.n641 VSS 0.228728f
C3741 VDD.n642 VSS 0.07686f
C3742 VDD.n643 VSS 0.114689f
C3743 VDD.n644 VSS 0.11402f
C3744 VDD.n645 VSS 0.041108f
C3745 VDD.n646 VSS 0.16955f
C3746 VDD.n647 VSS 0.169009f
C3747 VDD.n648 VSS 0.090794f
C3748 VDD.n649 VSS 0.114961f
C3749 VDD.n650 VSS 0.077132f
C3750 VDD.n651 VSS 0.299991f
C3751 VDD.n652 VSS 0.228728f
C3752 VDD.n653 VSS 0.07686f
C3753 VDD.n654 VSS 0.114689f
C3754 VDD.n655 VSS 0.11402f
C3755 VDD.n656 VSS 0.041108f
C3756 VDD.n657 VSS 0.16955f
C3757 VDD.n658 VSS 0.169009f
C3758 VDD.n659 VSS 0.090794f
C3759 VDD.n660 VSS 0.114961f
C3760 VDD.n661 VSS 0.077132f
C3761 VDD.n662 VSS 0.299991f
C3762 VDD.n663 VSS 0.228728f
C3763 VDD.n664 VSS 0.07686f
C3764 VDD.n665 VSS 0.114689f
C3765 VDD.n666 VSS 0.11402f
C3766 VDD.n667 VSS 0.041108f
C3767 VDD.n668 VSS 0.16955f
C3768 VDD.n669 VSS 0.169009f
C3769 VDD.n670 VSS 0.090794f
C3770 VDD.n671 VSS 0.114961f
C3771 VDD.n672 VSS 0.077132f
C3772 VDD.n673 VSS 0.299991f
C3773 VDD.n674 VSS 0.228728f
C3774 VDD.n675 VSS 0.07686f
C3775 VDD.n676 VSS 0.114689f
C3776 VDD.n677 VSS 0.11402f
C3777 VDD.n678 VSS 0.041108f
C3778 VDD.n679 VSS 0.16955f
C3779 VDD.n680 VSS 0.169009f
C3780 VDD.n681 VSS 0.090794f
C3781 VDD.n682 VSS 0.114961f
C3782 VDD.n683 VSS 0.077132f
C3783 VDD.n684 VSS 0.299991f
C3784 VDD.n685 VSS 0.228728f
C3785 VDD.n686 VSS 0.07686f
C3786 VDD.n687 VSS 0.114689f
C3787 VDD.n688 VSS 0.11402f
C3788 VDD.n689 VSS 0.041108f
C3789 VDD.n690 VSS 0.16955f
C3790 VDD.n691 VSS 0.169009f
C3791 VDD.n692 VSS 0.090794f
C3792 VDD.n693 VSS 0.114961f
C3793 VDD.n694 VSS 0.077132f
C3794 VDD.n695 VSS 0.299991f
C3795 VDD.n696 VSS 0.228728f
C3796 VDD.n697 VSS 0.07686f
C3797 VDD.n698 VSS 0.114689f
C3798 VDD.n699 VSS 0.11402f
C3799 VDD.n700 VSS 0.041108f
C3800 VDD.n701 VSS 0.16955f
C3801 VDD.n702 VSS 0.169009f
C3802 VDD.n703 VSS 0.090794f
C3803 VDD.n704 VSS 0.114961f
C3804 VDD.n705 VSS 0.077132f
C3805 VDD.n706 VSS 0.299991f
C3806 VDD.n707 VSS 0.228728f
C3807 VDD.n708 VSS 0.07686f
C3808 VDD.n709 VSS 0.114689f
C3809 VDD.n710 VSS 0.11402f
C3810 VDD.n711 VSS 0.041108f
C3811 VDD.n712 VSS 0.16955f
C3812 VDD.n713 VSS 0.169009f
C3813 VDD.n714 VSS 0.113512f
C3814 VDD.n715 VSS 0.114689f
C3815 VDD.t9 VSS 0.019607f
C3816 VDD.t65 VSS 0.019607f
C3817 VDD.n716 VSS 0.041911f
C3818 VDD.t269 VSS 0.019607f
C3819 VDD.t451 VSS 0.019607f
C3820 VDD.n717 VSS 0.041911f
C3821 VDD.t480 VSS 0.019607f
C3822 VDD.t289 VSS 0.019607f
C3823 VDD.n718 VSS 0.041911f
C3824 VDD.n719 VSS 0.16955f
C3825 VDD.n720 VSS 0.138239f
C3826 VDD.n721 VSS 0.132598f
C3827 VDD.n722 VSS 0.07686f
C3828 VDD.n723 VSS 0.114689f
C3829 VDD.t255 VSS 0.019607f
C3830 VDD.t217 VSS 0.019607f
C3831 VDD.n724 VSS 0.041911f
C3832 VDD.t443 VSS 0.019607f
C3833 VDD.t99 VSS 0.019607f
C3834 VDD.n725 VSS 0.041911f
C3835 VDD.t97 VSS 0.019607f
C3836 VDD.t259 VSS 0.019607f
C3837 VDD.n726 VSS 0.041911f
C3838 VDD.n727 VSS 0.16955f
C3839 VDD.n728 VSS 0.138239f
C3840 VDD.n729 VSS 0.132598f
C3841 VDD.n730 VSS 0.07686f
C3842 VDD.n731 VSS 0.114689f
C3843 VDD.t325 VSS 0.019607f
C3844 VDD.t327 VSS 0.019607f
C3845 VDD.n732 VSS 0.041911f
C3846 VDD.t130 VSS 0.019607f
C3847 VDD.t355 VSS 0.019607f
C3848 VDD.n733 VSS 0.041911f
C3849 VDD.t79 VSS 0.019607f
C3850 VDD.t497 VSS 0.019607f
C3851 VDD.n734 VSS 0.041911f
C3852 VDD.n735 VSS 0.16955f
C3853 VDD.n736 VSS 0.138239f
C3854 VDD.n737 VSS 0.132598f
C3855 VDD.n738 VSS 0.07686f
C3856 VDD.n739 VSS 0.114689f
C3857 VDD.t382 VSS 0.019607f
C3858 VDD.t380 VSS 0.019607f
C3859 VDD.n740 VSS 0.041911f
C3860 VDD.t347 VSS 0.019607f
C3861 VDD.t12 VSS 0.019607f
C3862 VDD.n741 VSS 0.041911f
C3863 VDD.t359 VSS 0.019607f
C3864 VDD.t414 VSS 0.019607f
C3865 VDD.n742 VSS 0.041911f
C3866 VDD.n743 VSS 0.16955f
C3867 VDD.n744 VSS 0.138239f
C3868 VDD.n745 VSS 0.132598f
C3869 VDD.n746 VSS 0.07686f
C3870 VDD.n747 VSS 0.114689f
C3871 VDD.t499 VSS 0.019607f
C3872 VDD.t253 VSS 0.019607f
C3873 VDD.n748 VSS 0.041911f
C3874 VDD.t501 VSS 0.019607f
C3875 VDD.t400 VSS 0.019607f
C3876 VDD.n749 VSS 0.041911f
C3877 VDD.t464 VSS 0.019607f
C3878 VDD.t339 VSS 0.019607f
C3879 VDD.n750 VSS 0.041911f
C3880 VDD.n751 VSS 0.16955f
C3881 VDD.n752 VSS 0.138239f
C3882 VDD.n753 VSS 0.132598f
C3883 VDD.n754 VSS 0.07686f
C3884 VDD.n755 VSS 0.114689f
C3885 VDD.t55 VSS 0.019607f
C3886 VDD.t386 VSS 0.019607f
C3887 VDD.n756 VSS 0.041911f
C3888 VDD.t126 VSS 0.019607f
C3889 VDD.t257 VSS 0.019607f
C3890 VDD.n757 VSS 0.041911f
C3891 VDD.t331 VSS 0.019607f
C3892 VDD.t293 VSS 0.019607f
C3893 VDD.n758 VSS 0.041911f
C3894 VDD.n759 VSS 0.16955f
C3895 VDD.n760 VSS 0.138239f
C3896 VDD.n761 VSS 0.132598f
C3897 VDD.n762 VSS 0.07686f
C3898 VDD.n763 VSS 0.114689f
C3899 VDD.t47 VSS 0.019607f
C3900 VDD.t378 VSS 0.019607f
C3901 VDD.n764 VSS 0.041911f
C3902 VDD.t449 VSS 0.019607f
C3903 VDD.t173 VSS 0.019607f
C3904 VDD.n765 VSS 0.041911f
C3905 VDD.t122 VSS 0.019607f
C3906 VDD.t95 VSS 0.019607f
C3907 VDD.n766 VSS 0.041911f
C3908 VDD.n767 VSS 0.16955f
C3909 VDD.n768 VSS 0.138239f
C3910 VDD.n769 VSS 0.132598f
C3911 VDD.n770 VSS 0.07686f
C3912 VDD.n771 VSS 0.114689f
C3913 VDD.t337 VSS 0.019607f
C3914 VDD.t437 VSS 0.019607f
C3915 VDD.n772 VSS 0.041911f
C3916 VDD.t184 VSS 0.019607f
C3917 VDD.t236 VSS 0.019607f
C3918 VDD.n773 VSS 0.041911f
C3919 VDD.t279 VSS 0.019607f
C3920 VDD.t283 VSS 0.019607f
C3921 VDD.n774 VSS 0.041911f
C3922 VDD.n775 VSS 0.16955f
C3923 VDD.n776 VSS 0.138239f
C3924 VDD.n777 VSS 0.132598f
C3925 VDD.n778 VSS 0.07686f
C3926 VDD.n779 VSS 0.114689f
C3927 VDD.t73 VSS 0.019607f
C3928 VDD.t57 VSS 0.019607f
C3929 VDD.n780 VSS 0.041911f
C3930 VDD.t118 VSS 0.019607f
C3931 VDD.t490 VSS 0.019607f
C3932 VDD.n781 VSS 0.041911f
C3933 VDD.t309 VSS 0.019607f
C3934 VDD.t311 VSS 0.019607f
C3935 VDD.n782 VSS 0.041911f
C3936 VDD.n783 VSS 0.16955f
C3937 VDD.n784 VSS 0.138239f
C3938 VDD.n785 VSS 0.132598f
C3939 VDD.n786 VSS 0.07686f
C3940 VDD.t410 VSS 0.019607f
C3941 VDD.t394 VSS 0.019607f
C3942 VDD.n787 VSS 0.041911f
C3943 VDD.n788 VSS 0.243627f
C3944 VDD.n789 VSS 0.12443f
C3945 VDD.n790 VSS 0.335724f
C3946 VDD.t409 VSS 0.300011f
C3947 VDD.t393 VSS 0.202292f
C3948 VDD.t308 VSS 0.202292f
C3949 VDD.t310 VSS 0.268957f
C3950 VDD.n791 VSS 0.100553f
C3951 VDD.n792 VSS 0.172408f
C3952 VDD.n793 VSS 0.228728f
C3953 VDD.t56 VSS 0.267808f
C3954 VDD.t72 VSS 0.202292f
C3955 VDD.t489 VSS 0.202292f
C3956 VDD.t117 VSS 0.264359f
C3957 VDD.n794 VSS 0.167811f
C3958 VDD.n795 VSS 0.11402f
C3959 VDD.n796 VSS 0.11402f
C3960 VDD.n797 VSS 0.041108f
C3961 VDD.n798 VSS 0.168684f
C3962 VDD.n799 VSS 0.169009f
C3963 VDD.n800 VSS 0.199189f
C3964 VDD.t281 VSS 0.019607f
C3965 VDD.t71 VSS 0.019607f
C3966 VDD.n801 VSS 0.041911f
C3967 VDD.n802 VSS 0.169009f
C3968 VDD.n803 VSS 0.199189f
C3969 VDD.n804 VSS 0.114961f
C3970 VDD.n805 VSS 0.335724f
C3971 VDD.t280 VSS 0.300011f
C3972 VDD.t70 VSS 0.202292f
C3973 VDD.t278 VSS 0.202292f
C3974 VDD.t282 VSS 0.268957f
C3975 VDD.n806 VSS 0.100553f
C3976 VDD.n807 VSS 0.172408f
C3977 VDD.n808 VSS 0.228728f
C3978 VDD.t436 VSS 0.267808f
C3979 VDD.t336 VSS 0.202292f
C3980 VDD.t235 VSS 0.202292f
C3981 VDD.t183 VSS 0.264359f
C3982 VDD.n809 VSS 0.167811f
C3983 VDD.n810 VSS 0.11402f
C3984 VDD.n811 VSS 0.11402f
C3985 VDD.n812 VSS 0.041108f
C3986 VDD.n813 VSS 0.168684f
C3987 VDD.n814 VSS 0.169009f
C3988 VDD.n815 VSS 0.199189f
C3989 VDD.t93 VSS 0.019607f
C3990 VDD.t63 VSS 0.019607f
C3991 VDD.n816 VSS 0.041911f
C3992 VDD.n817 VSS 0.169009f
C3993 VDD.n818 VSS 0.199189f
C3994 VDD.n819 VSS 0.114961f
C3995 VDD.n820 VSS 0.335724f
C3996 VDD.t92 VSS 0.300011f
C3997 VDD.t62 VSS 0.202292f
C3998 VDD.t121 VSS 0.202292f
C3999 VDD.t94 VSS 0.268957f
C4000 VDD.n821 VSS 0.100553f
C4001 VDD.n822 VSS 0.172408f
C4002 VDD.n823 VSS 0.228728f
C4003 VDD.t377 VSS 0.267808f
C4004 VDD.t46 VSS 0.202292f
C4005 VDD.t172 VSS 0.202292f
C4006 VDD.t448 VSS 0.264359f
C4007 VDD.n824 VSS 0.167811f
C4008 VDD.n825 VSS 0.11402f
C4009 VDD.n826 VSS 0.11402f
C4010 VDD.n827 VSS 0.041108f
C4011 VDD.n828 VSS 0.168684f
C4012 VDD.n829 VSS 0.169009f
C4013 VDD.n830 VSS 0.199189f
C4014 VDD.t299 VSS 0.019607f
C4015 VDD.t112 VSS 0.019607f
C4016 VDD.n831 VSS 0.041911f
C4017 VDD.n832 VSS 0.169009f
C4018 VDD.n833 VSS 0.199189f
C4019 VDD.n834 VSS 0.114961f
C4020 VDD.n835 VSS 0.335724f
C4021 VDD.t298 VSS 0.300011f
C4022 VDD.t111 VSS 0.202292f
C4023 VDD.t330 VSS 0.202292f
C4024 VDD.t292 VSS 0.268957f
C4025 VDD.n836 VSS 0.100553f
C4026 VDD.n837 VSS 0.172408f
C4027 VDD.n838 VSS 0.228728f
C4028 VDD.t385 VSS 0.267808f
C4029 VDD.t54 VSS 0.202292f
C4030 VDD.t256 VSS 0.202292f
C4031 VDD.t125 VSS 0.264359f
C4032 VDD.n839 VSS 0.167811f
C4033 VDD.n840 VSS 0.11402f
C4034 VDD.n841 VSS 0.11402f
C4035 VDD.n842 VSS 0.041108f
C4036 VDD.n843 VSS 0.168684f
C4037 VDD.n844 VSS 0.169009f
C4038 VDD.n845 VSS 0.199189f
C4039 VDD.t474 VSS 0.019607f
C4040 VDD.t372 VSS 0.019607f
C4041 VDD.n846 VSS 0.041911f
C4042 VDD.n847 VSS 0.169009f
C4043 VDD.n848 VSS 0.199189f
C4044 VDD.n849 VSS 0.114961f
C4045 VDD.n850 VSS 0.335724f
C4046 VDD.t473 VSS 0.300011f
C4047 VDD.t371 VSS 0.202292f
C4048 VDD.t463 VSS 0.202292f
C4049 VDD.t338 VSS 0.268957f
C4050 VDD.n851 VSS 0.100553f
C4051 VDD.n852 VSS 0.172408f
C4052 VDD.n853 VSS 0.228728f
C4053 VDD.t252 VSS 0.267808f
C4054 VDD.t498 VSS 0.202292f
C4055 VDD.t399 VSS 0.202292f
C4056 VDD.t500 VSS 0.264359f
C4057 VDD.n854 VSS 0.167811f
C4058 VDD.n855 VSS 0.11402f
C4059 VDD.n856 VSS 0.11402f
C4060 VDD.n857 VSS 0.041108f
C4061 VDD.n858 VSS 0.168684f
C4062 VDD.n859 VSS 0.169009f
C4063 VDD.n860 VSS 0.199189f
C4064 VDD.t482 VSS 0.019607f
C4065 VDD.t412 VSS 0.019607f
C4066 VDD.n861 VSS 0.041911f
C4067 VDD.n862 VSS 0.169009f
C4068 VDD.n863 VSS 0.199189f
C4069 VDD.n864 VSS 0.114961f
C4070 VDD.n865 VSS 0.335724f
C4071 VDD.t481 VSS 0.300011f
C4072 VDD.t411 VSS 0.202292f
C4073 VDD.t358 VSS 0.202292f
C4074 VDD.t413 VSS 0.268957f
C4075 VDD.n866 VSS 0.100553f
C4076 VDD.n867 VSS 0.172408f
C4077 VDD.n868 VSS 0.228728f
C4078 VDD.t379 VSS 0.267808f
C4079 VDD.t381 VSS 0.202292f
C4080 VDD.t11 VSS 0.202292f
C4081 VDD.t346 VSS 0.264359f
C4082 VDD.n869 VSS 0.167811f
C4083 VDD.n870 VSS 0.11402f
C4084 VDD.n871 VSS 0.11402f
C4085 VDD.n872 VSS 0.041108f
C4086 VDD.n873 VSS 0.168684f
C4087 VDD.n874 VSS 0.169009f
C4088 VDD.n875 VSS 0.199189f
C4089 VDD.t182 VSS 0.019607f
C4090 VDD.t77 VSS 0.019607f
C4091 VDD.n876 VSS 0.041911f
C4092 VDD.n877 VSS 0.169009f
C4093 VDD.n878 VSS 0.199189f
C4094 VDD.n879 VSS 0.114961f
C4095 VDD.n880 VSS 0.335724f
C4096 VDD.t181 VSS 0.300011f
C4097 VDD.t76 VSS 0.202292f
C4098 VDD.t78 VSS 0.202292f
C4099 VDD.t496 VSS 0.268957f
C4100 VDD.n881 VSS 0.100553f
C4101 VDD.n882 VSS 0.172408f
C4102 VDD.n883 VSS 0.228728f
C4103 VDD.t326 VSS 0.267808f
C4104 VDD.t324 VSS 0.202292f
C4105 VDD.t354 VSS 0.202292f
C4106 VDD.t129 VSS 0.264359f
C4107 VDD.n884 VSS 0.167811f
C4108 VDD.n885 VSS 0.11402f
C4109 VDD.n886 VSS 0.11402f
C4110 VDD.n887 VSS 0.041108f
C4111 VDD.n888 VSS 0.168684f
C4112 VDD.n889 VSS 0.169009f
C4113 VDD.n890 VSS 0.199189f
C4114 VDD.t370 VSS 0.019607f
C4115 VDD.t186 VSS 0.019607f
C4116 VDD.n891 VSS 0.041911f
C4117 VDD.n892 VSS 0.169009f
C4118 VDD.n893 VSS 0.199189f
C4119 VDD.n894 VSS 0.114961f
C4120 VDD.n895 VSS 0.335724f
C4121 VDD.t369 VSS 0.300011f
C4122 VDD.t185 VSS 0.202292f
C4123 VDD.t96 VSS 0.202292f
C4124 VDD.t258 VSS 0.268957f
C4125 VDD.n896 VSS 0.100553f
C4126 VDD.n897 VSS 0.172408f
C4127 VDD.n898 VSS 0.228728f
C4128 VDD.t216 VSS 0.267808f
C4129 VDD.t254 VSS 0.202292f
C4130 VDD.t98 VSS 0.202292f
C4131 VDD.t442 VSS 0.264359f
C4132 VDD.n899 VSS 0.167811f
C4133 VDD.n900 VSS 0.11402f
C4134 VDD.n901 VSS 0.11402f
C4135 VDD.n902 VSS 0.041108f
C4136 VDD.n903 VSS 0.168684f
C4137 VDD.n904 VSS 0.169009f
C4138 VDD.n905 VSS 0.199189f
C4139 VDD.t211 VSS 0.019607f
C4140 VDD.t295 VSS 0.019607f
C4141 VDD.n906 VSS 0.041911f
C4142 VDD.n907 VSS 0.169009f
C4143 VDD.n908 VSS 0.199189f
C4144 VDD.n909 VSS 0.114961f
C4145 VDD.n910 VSS 0.335724f
C4146 VDD.t210 VSS 0.300011f
C4147 VDD.t294 VSS 0.202292f
C4148 VDD.t479 VSS 0.202292f
C4149 VDD.t288 VSS 0.268957f
C4150 VDD.n911 VSS 0.100553f
C4151 VDD.n912 VSS 0.172408f
C4152 VDD.n913 VSS 0.228728f
C4153 VDD.t64 VSS 0.267808f
C4154 VDD.t8 VSS 0.202292f
C4155 VDD.t450 VSS 0.202292f
C4156 VDD.t268 VSS 0.264359f
C4157 VDD.n914 VSS 0.167811f
C4158 VDD.n915 VSS 0.11402f
C4159 VDD.n916 VSS 0.11402f
C4160 VDD.n917 VSS 0.041108f
C4161 VDD.n918 VSS 0.168684f
C4162 VDD.n919 VSS 0.169009f
C4163 VDD.n920 VSS 0.132767f
C4164 VDD.n921 VSS 0.121664f
C4165 VDD.n922 VSS 0.470659f
C4166 VDD.n923 VSS 0.793242f
C4167 VDD.n924 VSS 0.085001f
C4168 VDD.n925 VSS 0.146538f
C4169 VDD.n926 VSS 0.387327f
C4170 VDD.t296 VSS 0.301845f
C4171 VDD.t260 VSS 0.190393f
C4172 VDD.t180 VSS 0.190393f
C4173 VDD.t189 VSS 0.249891f
C4174 VDD.n927 VSS 0.156858f
C4175 VDD.n928 VSS 0.043203f
C4176 VDD.n929 VSS 0.159021f
C4177 VDD.t233 VSS 0.252054f
C4178 VDD.t251 VSS 0.190393f
C4179 VDD.t290 VSS 0.190393f
C4180 VDD.t348 VSS 0.296651f
C4181 VDD.n930 VSS 0.383723f
C4182 VDD.n931 VSS 0.100844f
C4183 VDD.n932 VSS 0.146538f
C4184 VDD.n933 VSS 0.129206f
C4185 VDD.n934 VSS 0.011609f
C4186 VDD.n935 VSS 0.170163f
C4187 VDD.n936 VSS 0.174348f
C4188 VDD.n937 VSS 0.137873f
C4189 VDD.n938 VSS 0.085001f
C4190 VDD.n939 VSS 0.146538f
C4191 VDD.n940 VSS 0.387327f
C4192 VDD.t342 VSS 0.301845f
C4193 VDD.t397 VSS 0.190393f
C4194 VDD.t494 VSS 0.190393f
C4195 VDD.t156 VSS 0.249891f
C4196 VDD.n941 VSS 0.156858f
C4197 VDD.n942 VSS 0.043203f
C4198 VDD.n943 VSS 0.159021f
C4199 VDD.t270 VSS 0.252054f
C4200 VDD.t10 VSS 0.190393f
C4201 VDD.t225 VSS 0.190393f
C4202 VDD.t135 VSS 0.296651f
C4203 VDD.n944 VSS 0.383723f
C4204 VDD.n945 VSS 0.100844f
C4205 VDD.n946 VSS 0.146538f
C4206 VDD.n947 VSS 0.129206f
C4207 VDD.n948 VSS 0.011609f
C4208 VDD.n949 VSS 0.170163f
C4209 VDD.n950 VSS 0.174348f
C4210 VDD.n951 VSS 0.137873f
C4211 VDD.n952 VSS 0.085001f
C4212 VDD.n953 VSS 0.146538f
C4213 VDD.n954 VSS 0.387327f
C4214 VDD.t444 VSS 0.301845f
C4215 VDD.t137 VSS 0.190393f
C4216 VDD.t248 VSS 0.190393f
C4217 VDD.t286 VSS 0.249891f
C4218 VDD.n955 VSS 0.156858f
C4219 VDD.n956 VSS 0.043203f
C4220 VDD.n957 VSS 0.159021f
C4221 VDD.t193 VSS 0.252054f
C4222 VDD.t149 VSS 0.190393f
C4223 VDD.t458 VSS 0.190393f
C4224 VDD.t274 VSS 0.296651f
C4225 VDD.n958 VSS 0.383723f
C4226 VDD.n959 VSS 0.100844f
C4227 VDD.n960 VSS 0.146538f
C4228 VDD.n961 VSS 0.129206f
C4229 VDD.n962 VSS 0.011609f
C4230 VDD.n963 VSS 0.170163f
C4231 VDD.n964 VSS 0.174348f
C4232 VDD.n965 VSS 0.137873f
C4233 VDD.n966 VSS 0.085001f
C4234 VDD.n967 VSS 0.146538f
C4235 VDD.n968 VSS 0.387327f
C4236 VDD.t0 VSS 0.301845f
C4237 VDD.t139 VSS 0.190393f
C4238 VDD.t224 VSS 0.190393f
C4239 VDD.t469 VSS 0.249891f
C4240 VDD.n969 VSS 0.156858f
C4241 VDD.n970 VSS 0.043203f
C4242 VDD.n971 VSS 0.159021f
C4243 VDD.t387 VSS 0.252054f
C4244 VDD.t239 VSS 0.190393f
C4245 VDD.t4 VSS 0.190393f
C4246 VDD.t141 VSS 0.296651f
C4247 VDD.n972 VSS 0.383723f
C4248 VDD.n973 VSS 0.100844f
C4249 VDD.n974 VSS 0.146538f
C4250 VDD.n975 VSS 0.129206f
C4251 VDD.n976 VSS 0.011609f
C4252 VDD.n977 VSS 0.170163f
C4253 VDD.n978 VSS 0.174348f
C4254 VDD.n979 VSS 0.137873f
C4255 VDD.n980 VSS 0.085001f
C4256 VDD.n981 VSS 0.146538f
C4257 VDD.n982 VSS 0.387327f
C4258 VDD.t419 VSS 0.301845f
C4259 VDD.t421 VSS 0.190393f
C4260 VDD.t491 VSS 0.190393f
C4261 VDD.t24 VSS 0.249891f
C4262 VDD.n983 VSS 0.156858f
C4263 VDD.n984 VSS 0.043203f
C4264 VDD.n985 VSS 0.159021f
C4265 VDD.t154 VSS 0.252054f
C4266 VDD.t433 VSS 0.190393f
C4267 VDD.t425 VSS 0.190393f
C4268 VDD.t427 VSS 0.296651f
C4269 VDD.n986 VSS 0.383723f
C4270 VDD.n987 VSS 0.100844f
C4271 VDD.n988 VSS 0.146538f
C4272 VDD.n989 VSS 0.129206f
C4273 VDD.n990 VSS 0.011609f
C4274 VDD.n991 VSS 0.170163f
C4275 VDD.n992 VSS 0.174348f
C4276 VDD.n993 VSS 0.137873f
C4277 VDD.n994 VSS 0.085001f
C4278 VDD.n995 VSS 0.146538f
C4279 VDD.n996 VSS 0.387327f
C4280 VDD.t328 VSS 0.301845f
C4281 VDD.t58 VSS 0.190393f
C4282 VDD.t462 VSS 0.190393f
C4283 VDD.t127 VSS 0.249891f
C4284 VDD.n997 VSS 0.156858f
C4285 VDD.n998 VSS 0.043203f
C4286 VDD.n999 VSS 0.159021f
C4287 VDD.t383 VSS 0.252054f
C4288 VDD.t110 VSS 0.190393f
C4289 VDD.t391 VSS 0.190393f
C4290 VDD.t389 VSS 0.296651f
C4291 VDD.n1000 VSS 0.383723f
C4292 VDD.n1001 VSS 0.100844f
C4293 VDD.n1002 VSS 0.146538f
C4294 VDD.n1003 VSS 0.129206f
C4295 VDD.n1004 VSS 0.011609f
C4296 VDD.n1005 VSS 0.170163f
C4297 VDD.n1006 VSS 0.174348f
C4298 VDD.n1007 VSS 0.137873f
C4299 VDD.n1008 VSS 0.085001f
C4300 VDD.n1009 VSS 0.146538f
C4301 VDD.n1010 VSS 0.387327f
C4302 VDD.t362 VSS 0.301845f
C4303 VDD.t438 VSS 0.190393f
C4304 VDD.t15 VSS 0.190393f
C4305 VDD.t82 VSS 0.249891f
C4306 VDD.n1011 VSS 0.156858f
C4307 VDD.n1012 VSS 0.043203f
C4308 VDD.n1013 VSS 0.159021f
C4309 VDD.t434 VSS 0.252054f
C4310 VDD.t368 VSS 0.190393f
C4311 VDD.t360 VSS 0.190393f
C4312 VDD.t366 VSS 0.296651f
C4313 VDD.n1014 VSS 0.383723f
C4314 VDD.n1015 VSS 0.100844f
C4315 VDD.n1016 VSS 0.146538f
C4316 VDD.n1017 VSS 0.129206f
C4317 VDD.n1018 VSS 0.011609f
C4318 VDD.n1019 VSS 0.170163f
C4319 VDD.n1020 VSS 0.174348f
C4320 VDD.n1021 VSS 0.137873f
C4321 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n0 VSS 1.0614f
C4322 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t6 VSS 0.096169f
C4323 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t5 VSS 0.041341f
C4324 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n1 VSS 0.116331f
C4325 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t1 VSS 0.054421f
C4326 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t2 VSS 0.054421f
C4327 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n2 VSS 0.114315f
C4328 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t0 VSS 0.202807f
C4329 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t3 VSS 0.200111f
C4330 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t10 VSS 0.087824f
C4331 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t7 VSS 0.040008f
C4332 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n3 VSS 0.097717f
C4333 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n4 VSS 0.382243f
C4334 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t4 VSS 0.107599f
C4335 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n5 VSS 0.139678f
C4336 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t8 VSS 0.082007f
C4337 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.t9 VSS 0.090862f
C4338 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n6 VSS 0.108213f
C4339 vernier_delay_line_0.saff_delay_unit_6/saff_2_0.sense_amplifier_0.out1.n7 VSS 1.24645f
.ends

