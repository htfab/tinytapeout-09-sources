magic
tech sky130A
magscale 1 2
timestamp 1731171178
<< nmos >>
rect -15 -200 15 200
<< ndiff >>
rect -73 188 -15 200
rect -73 -188 -61 188
rect -27 -188 -15 188
rect -73 -200 -15 -188
rect 15 188 73 200
rect 15 -188 27 188
rect 61 -188 73 188
rect 15 -200 73 -188
<< ndiffc >>
rect -61 -188 -27 188
rect 27 -188 61 188
<< poly >>
rect -15 200 15 226
rect -15 -226 15 -200
<< locali >>
rect -61 188 -27 204
rect -61 -204 -27 -188
rect 27 188 61 204
rect 27 -204 61 -188
<< viali >>
rect -61 -188 -27 188
rect 27 -188 61 188
<< metal1 >>
rect -67 188 -21 200
rect -67 -188 -61 188
rect -27 -188 -21 188
rect -67 -200 -21 -188
rect 21 188 67 200
rect 21 -188 27 188
rect 61 -188 67 188
rect 21 -200 67 -188
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
