magic
tech sky130A
timestamp 1730750158
use inverter_3_1  inverter_3_1_0
timestamp 1730749971
transform 1 0 2 0 1 110
box 15 -98 214 543
use inverter_3_1  inverter_3_1_2
timestamp 1730749971
transform 1 0 147 0 1 110
box 15 -98 214 543
use inverter_3_1  inverter_3_1_3
timestamp 1730749971
transform 1 0 292 0 1 110
box 15 -98 214 543
use inverter_3_1  inverter_3_1_4
timestamp 1730749971
transform 1 0 437 0 1 110
box 15 -98 214 543
<< end >>
