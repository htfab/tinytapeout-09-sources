magic
tech sky130A
magscale 1 2
timestamp 1730882523
<< pwell >>
rect -201 -652 201 652
<< psubdiff >>
rect -165 582 -69 616
rect 69 582 165 616
rect -165 520 -131 582
rect 131 520 165 582
rect -165 -582 -131 -520
rect 131 -582 165 -520
rect -165 -616 -69 -582
rect 69 -616 165 -582
<< psubdiffcont >>
rect -69 582 69 616
rect -165 -520 -131 520
rect 131 -520 165 520
rect -69 -616 69 -582
<< xpolycontact >>
rect -35 54 35 486
rect -35 -486 35 -54
<< xpolyres >>
rect -35 -54 35 54
<< locali >>
rect -165 582 -69 616
rect 69 582 165 616
rect -165 520 -131 582
rect 131 520 165 582
rect -165 -582 -131 -520
rect 131 -582 165 -520
rect -165 -616 -69 -582
rect 69 -616 165 -582
<< viali >>
rect -19 71 19 468
rect -19 -468 19 -71
<< metal1 >>
rect -25 468 25 480
rect -25 71 -19 468
rect 19 71 25 468
rect -25 59 25 71
rect -25 -71 25 -59
rect -25 -468 -19 -71
rect 19 -468 25 -71
rect -25 -480 25 -468
<< properties >>
string FIXED_BBOX -148 -599 148 599
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.7 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
