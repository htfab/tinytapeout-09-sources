*SWTCH_INV_SKY130NM/SWTCH_INV
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/SWTCH_INV_lpe.spi
#else
.include ../../../work/xsch/SWTCH_INV.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VDD  VDD  GND  pwl 0 0 1p {AVDD}

VIN  IN   GND  pwl 0 0 1n 0 2n {AVDD} 5n {AVDD} 6n 0

Rload OUT GND 100k

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD GND IN OUT SWTCH_INV

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.probe v(VDD) v(GND) v(IN) v(OUT)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 10n 1p
write
quit
#endif

.endc

.end
