** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/input_stage.sch
.subckt input_stage in en t0 t1 t2 t3 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B t0:I t1:I t2:I t3:I en:I
x1 en in net1 VDD VSS nand_gate
x2 net1 net2 VDD VSS inverter_2
x3 net2 t0 t1 net3 VDD VSS fine_delay
x4 net3 t2 t3 out VDD VSS fine_delay
.ends

* expanding   symbol:  nand_gate.sym # of pins=5
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/nand_gate.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/nand_gate.sch
.subckt nand_gate a b out VDD VSS
*.PININFO VDD:B a:I out:O VSS:B b:I
XM7 out a net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM1 out a VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net1 b VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 out b VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
.ends


* expanding   symbol:  inverter_2.sym # of pins=4
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/inverter_2.sch
.subckt inverter_2 in out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B
XM1 out in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 out in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends


* expanding   symbol:  fine_delay.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/fine_delay.sym
** sch_path: /home/ttuser/Documents/tt09-analog-tdc/xschem/fine_delay.sch
.subckt fine_delay in t0 t1 out VDD VSS
*.PININFO VDD:B in:I out:O VSS:B t0:I t1:I
XM1 net1 in VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM2 net3 in VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 net3 t1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM8 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM9 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM10 net2 in net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM11 net2 t0 net3 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=2 nf=1 m=1
XM3 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net1 in net2 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends

.end
