* NGSPICE file created from nand_gate_parax.ext - technology: sky130A

.subckt nand_gate_parax a b out VDD VSS
X0 out.t0 a.t0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X1 VDD.t3 b.t0 out.t2 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X2 VSS.t2 b.t1 a_124_n546# VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.15
X3 a_124_n546# a.t1 out.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.15
R0 a.n0 a.t0 564.04
R1 a.n0 a.t1 511.623
R2 a a.n0 161.375
R3 VDD.n6 VDD.n3 1348.04
R4 VDD.n6 VDD.n4 1348.04
R5 VDD.t0 VDD.n4 181.043
R6 VDD.t2 VDD.n3 176.736
R7 VDD.n7 VDD.n0 143.792
R8 VDD.n7 VDD.n2 143.792
R9 VDD.n9 VDD.t1 84.7879
R10 VDD.n1 VDD.t3 84.7879
R11 VDD.n5 VDD.t2 49.547
R12 VDD.n5 VDD.t0 45.2386
R13 VDD.n4 VDD.n0 20.5561
R14 VDD.n3 VDD.n2 20.5561
R15 VDD.n7 VDD.n6 18.5005
R16 VDD.n6 VDD.n5 18.5005
R17 VDD.n2 VDD.n1 2.16438
R18 VDD.n10 VDD.n0 2.0406
R19 VDD.n8 VDD.n7 1.8605
R20 VDD.n10 VDD.n9 0.129176
R21 VDD.n8 VDD.n1 0.110794
R22 VDD.n9 VDD.n8 0.105892
R23 VDD VDD.n10 0.0666765
R24 out.n1 out.n0 75.7065
R25 out.n1 out.t1 42.0134
R26 out.n0 out.t2 9.52217
R27 out.n0 out.t0 9.52217
R28 out out.n1 0.063
R29 b.n0 b.t0 618.668
R30 b.n0 b.t1 456.997
R31 b b.n0 161.333
R32 VSS.n6 VSS.n4 1707.33
R33 VSS.n6 VSS.n3 1707.33
R34 VSS.t1 VSS.n3 1000.06
R35 VSS.t0 VSS.n4 1000.06
R36 VSS.n5 VSS.t1 275.784
R37 VSS.n5 VSS.t0 275.784
R38 VSS.n7 VSS.n2 110.933
R39 VSS.n7 VSS.n0 110.933
R40 VSS.n3 VSS.n2 97.5005
R41 VSS.n4 VSS.n0 97.5005
R42 VSS.n7 VSS.n6 58.5005
R43 VSS.n6 VSS.n5 58.5005
R44 VSS.n1 VSS.t2 42.0841
R45 VSS.n2 VSS.n1 2.27599
R46 VSS.n9 VSS.n0 2.1305
R47 VSS.n8 VSS.n7 1.8605
R48 VSS.n9 VSS.n8 0.230892
R49 VSS.n8 VSS.n1 0.108343
R50 VSS VSS.n9 0.0728039
C0 VDD a_124_n546# 7.57e-19
C1 out a 0.114267f
C2 b a 0.078266f
C3 a a_124_n546# 0.009499f
C4 a VDD 0.135896f
C5 b out 0.050326f
C6 out a_124_n546# 0.355343f
C7 b a_124_n546# 0.009499f
C8 out VDD 1.0058f
C9 b VDD 0.116645f
C10 out VSS 0.429217f
C11 b VSS 0.249864f
C12 a VSS 0.197231f
C13 VDD VSS 2.21616f
C14 a_124_n546# VSS 0.371906f
.ends

