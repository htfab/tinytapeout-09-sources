magic
tech sky130A
magscale 1 2
timestamp 1731136808
<< nwell >>
rect 720 1352 1458 1570
rect 720 628 808 1352
rect 1290 628 1458 1352
<< pwell >>
rect 720 22 1458 628
<< psubdiff >>
rect 756 450 790 474
rect 1308 450 1342 474
rect 756 22 790 152
rect 1308 22 1342 152
<< nsubdiff >>
rect 756 1404 790 1534
rect 1308 1404 1342 1534
rect 756 686 790 710
rect 1308 686 1342 710
<< psubdiffcont >>
rect 756 152 790 450
rect 1308 152 1342 450
rect 790 22 1308 118
<< nsubdiffcont >>
rect 790 1438 1308 1534
rect 756 710 790 1404
rect 1308 710 1342 1404
<< poly >>
rect 970 1392 1044 1404
rect 970 1358 990 1392
rect 1024 1358 1044 1392
rect 970 1346 1044 1358
rect 902 1316 1108 1346
rect 1166 620 1196 664
rect 1088 608 1196 620
rect 1088 574 1108 608
rect 1142 574 1196 608
rect 1088 562 1196 574
rect 1166 496 1196 562
rect 902 214 1108 244
rect 968 202 1042 214
rect 968 168 988 202
rect 1022 168 1042 202
rect 968 156 1042 168
<< polycont >>
rect 990 1358 1024 1392
rect 1108 574 1142 608
rect 988 168 1022 202
<< locali >>
rect 756 1404 790 1534
rect 1308 1404 1342 1534
rect 970 1392 1044 1404
rect 970 1358 990 1392
rect 1024 1358 1044 1392
rect 970 1346 1044 1358
rect 756 686 790 710
rect 1308 686 1342 710
rect 1088 608 1162 620
rect 1088 574 1108 608
rect 1142 574 1162 608
rect 1088 562 1162 574
rect 756 450 790 474
rect 1308 450 1342 474
rect 968 202 1042 214
rect 968 168 988 202
rect 1022 168 1042 202
rect 968 156 1042 168
rect 756 22 790 152
rect 1308 22 1342 152
<< viali >>
rect 790 1444 1308 1528
rect 756 710 790 1404
rect 990 1358 1024 1392
rect 1308 710 1342 1404
rect 1108 574 1142 608
rect 756 152 790 450
rect 988 168 1022 202
rect 1308 152 1342 450
rect 790 28 1308 112
<< metal1 >>
rect 720 1528 1458 1534
rect 720 1444 790 1528
rect 1308 1444 1458 1528
rect 720 1438 1458 1444
rect 750 1404 796 1438
rect 750 710 756 1404
rect 790 710 796 1404
rect 850 1290 896 1438
rect 970 1406 1044 1410
rect 970 1344 976 1406
rect 1038 1344 1044 1406
rect 970 1340 1044 1344
rect 1302 1404 1348 1438
rect 930 1284 992 1290
rect 930 1192 934 1284
rect 988 1192 992 1284
rect 930 1186 992 1192
rect 1106 1284 1168 1290
rect 1106 1192 1110 1284
rect 1164 1192 1168 1284
rect 1106 1186 1168 1192
rect 750 686 796 710
rect 842 788 904 794
rect 842 696 846 788
rect 900 696 904 788
rect 842 690 904 696
rect 1018 788 1080 794
rect 1018 696 1022 788
rect 1076 696 1080 788
rect 1018 690 1080 696
rect 1302 710 1308 1404
rect 1342 710 1348 1404
rect 930 608 1162 620
rect 930 574 1108 608
rect 1142 574 1162 608
rect 930 562 1162 574
rect 1202 608 1248 690
rect 1302 686 1348 710
rect 1202 550 1458 608
rect 750 450 796 474
rect 1202 470 1248 550
rect 750 152 756 450
rect 790 152 796 450
rect 842 464 904 470
rect 842 402 846 464
rect 900 402 904 464
rect 842 396 904 402
rect 1018 464 1080 470
rect 1018 402 1022 464
rect 1076 402 1080 464
rect 1018 396 1080 402
rect 1302 450 1348 474
rect 930 338 992 344
rect 930 276 934 338
rect 988 276 992 338
rect 930 270 992 276
rect 1106 338 1168 344
rect 1106 276 1110 338
rect 1164 276 1168 338
rect 1106 270 1168 276
rect 750 118 796 152
rect 850 118 896 270
rect 968 216 1042 220
rect 968 154 974 216
rect 1036 154 1042 216
rect 968 150 1042 154
rect 1302 152 1308 450
rect 1342 152 1348 450
rect 1302 118 1348 152
rect 720 112 1458 118
rect 720 28 790 112
rect 1308 28 1458 112
rect 720 22 1458 28
<< via1 >>
rect 976 1392 1038 1406
rect 976 1358 990 1392
rect 990 1358 1024 1392
rect 1024 1358 1038 1392
rect 976 1344 1038 1358
rect 934 1192 988 1284
rect 1110 1192 1164 1284
rect 846 696 900 788
rect 1022 696 1076 788
rect 846 402 900 464
rect 1022 402 1076 464
rect 934 276 988 338
rect 1110 276 1164 338
rect 974 202 1036 216
rect 974 168 988 202
rect 988 168 1022 202
rect 1022 168 1036 202
rect 974 154 1036 168
<< metal2 >>
rect 970 1406 1044 1638
rect 970 1344 976 1406
rect 1038 1344 1044 1406
rect 970 1340 1044 1344
rect 930 1284 1168 1290
rect 930 1192 934 1284
rect 988 1192 1110 1284
rect 1164 1192 1168 1284
rect 930 1186 1168 1192
rect 842 788 1080 794
rect 842 696 846 788
rect 900 696 1022 788
rect 1076 696 1080 788
rect 842 690 1080 696
rect 842 464 1080 470
rect 842 402 846 464
rect 900 402 1022 464
rect 1076 402 1080 464
rect 842 396 1080 402
rect 930 338 1168 344
rect 930 276 934 338
rect 988 276 1110 338
rect 1164 276 1168 338
rect 930 270 1168 276
rect 1384 220 1454 1638
rect 968 216 1454 220
rect 968 154 974 216
rect 1036 154 1454 216
rect 968 150 1454 154
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1730191042
transform 1 0 917 0 1 370
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1730191042
transform 1 0 1005 0 1 370
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1730191042
transform 1 0 1093 0 1 370
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1730191042
transform 1 0 1181 0 1 370
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 917 0 1 990
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_1
timestamp 1730191042
transform 1 0 1005 0 1 990
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_2
timestamp 1730191042
transform 1 0 1093 0 1 990
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_3
timestamp 1730191042
transform 1 0 1181 0 1 990
box -109 -362 109 362
<< labels >>
rlabel metal1 930 562 988 620 0 in
port 1 nsew
rlabel metal2 1384 1580 1442 1638 0 en
port 2 nsew
rlabel metal2 970 1580 1028 1638 0 nen
port 3 nsew
rlabel metal1 1300 550 1358 608 0 out
port 4 nsew
rlabel metal1 720 1476 778 1534 0 VDD
port 5 nsew
rlabel metal1 720 60 778 118 0 VSS
port 6 nsew
<< end >>
