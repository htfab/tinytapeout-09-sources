magic
tech sky130A
magscale 1 2
timestamp 1730306345
<< error_p >>
rect -35 1070 35 1072
rect -35 34 35 36
rect -35 -1002 35 -1000
<< pwell >>
rect -201 -1668 201 1668
<< psubdiff >>
rect -165 1598 -69 1632
rect 69 1598 165 1632
rect -165 1536 -131 1598
rect 131 1536 165 1598
rect -165 -1598 -131 -1536
rect 131 -1598 165 -1536
rect -165 -1632 -69 -1598
rect 69 -1632 165 -1598
<< psubdiffcont >>
rect -69 1598 69 1632
rect -165 -1536 -131 1536
rect 131 -1536 165 1536
rect -69 -1632 69 -1598
<< xpolycontact >>
rect -35 1070 35 1502
rect -35 570 35 1002
rect -35 34 35 466
rect -35 -466 35 -34
rect -35 -1002 35 -570
rect -35 -1502 35 -1070
<< xpolyres >>
rect -35 1002 35 1070
rect -35 -34 35 34
rect -35 -1070 35 -1002
<< locali >>
rect -165 1598 -69 1632
rect 69 1598 165 1632
rect -165 1536 -131 1598
rect 131 1536 165 1598
rect -165 -1598 -131 -1536
rect 131 -1598 165 -1536
rect -165 -1632 -69 -1598
rect 69 -1632 165 -1598
<< viali >>
rect -19 1087 19 1484
rect -19 588 19 985
rect -19 51 19 448
rect -19 -448 19 -51
rect -19 -985 19 -588
rect -19 -1484 19 -1087
<< metal1 >>
rect -25 1484 25 1496
rect -25 1087 -19 1484
rect 19 1087 25 1484
rect -25 1075 25 1087
rect -25 985 25 997
rect -25 588 -19 985
rect 19 588 25 985
rect -25 576 25 588
rect -25 448 25 460
rect -25 51 -19 448
rect 19 51 25 448
rect -25 39 25 51
rect -25 -51 25 -39
rect -25 -448 -19 -51
rect 19 -448 25 -51
rect -25 -460 25 -448
rect -25 -588 25 -576
rect -25 -985 -19 -588
rect 19 -985 25 -588
rect -25 -997 25 -985
rect -25 -1087 25 -1075
rect -25 -1484 -19 -1087
rect 19 -1484 25 -1087
rect -25 -1496 25 -1484
<< properties >>
string FIXED_BBOX -148 -1615 148 1615
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.50 m 3 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
