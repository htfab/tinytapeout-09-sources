magic
tech sky130A
timestamp 1731256823
<< nwell >>
rect 334 2422 470 2558
<< pwell >>
rect 334 2558 470 2664
<< nmos >>
rect 410 2604 425 2646
<< pmoshvt >>
rect 410 2440 425 2540
<< ndiff >>
rect 380 2642 410 2646
rect 380 2608 387 2642
rect 404 2608 410 2642
rect 380 2604 410 2608
rect 425 2634 452 2646
rect 425 2616 431 2634
rect 448 2616 452 2634
rect 425 2604 452 2616
<< pdiff >>
rect 381 2536 410 2540
rect 381 2444 387 2536
rect 404 2444 410 2536
rect 381 2440 410 2444
rect 425 2528 452 2540
rect 425 2452 431 2528
rect 448 2452 452 2528
rect 425 2440 452 2452
<< ndiffc >>
rect 387 2608 404 2642
rect 431 2616 448 2634
<< pdiffc >>
rect 387 2444 404 2536
rect 431 2452 448 2528
<< psubdiff >>
rect 351 2634 380 2646
rect 351 2616 353 2634
rect 370 2616 380 2634
rect 351 2604 380 2616
<< nsubdiff >>
rect 352 2528 381 2540
rect 352 2452 353 2528
rect 370 2452 381 2528
rect 352 2440 381 2452
<< psubdiffcont >>
rect 353 2616 370 2634
<< nsubdiffcont >>
rect 353 2452 370 2528
<< poly >>
rect 410 2646 425 2659
rect 410 2586 425 2604
rect 392 2581 425 2586
rect 392 2564 400 2581
rect 417 2564 425 2581
rect 392 2559 425 2564
rect 410 2540 425 2559
rect 410 2427 425 2440
<< polycont >>
rect 400 2564 417 2581
<< locali >>
rect 345 2636 387 2642
rect 345 2614 348 2636
rect 345 2608 387 2614
rect 404 2608 412 2642
rect 431 2639 448 2642
rect 431 2608 448 2611
rect 417 2564 425 2581
rect 345 2530 387 2536
rect 345 2450 348 2530
rect 345 2444 387 2450
rect 404 2444 412 2536
rect 431 2533 448 2536
rect 431 2444 448 2447
<< viali >>
rect 348 2634 387 2636
rect 348 2616 353 2634
rect 353 2616 370 2634
rect 370 2616 387 2634
rect 348 2614 387 2616
rect 387 2614 402 2636
rect 431 2634 448 2639
rect 431 2616 448 2634
rect 431 2611 448 2616
rect 388 2564 400 2581
rect 400 2564 405 2581
rect 348 2528 387 2530
rect 348 2452 353 2528
rect 353 2452 370 2528
rect 370 2452 387 2528
rect 348 2450 387 2452
rect 387 2450 402 2530
rect 431 2528 448 2533
rect 431 2452 448 2528
rect 431 2447 448 2452
<< metal1 >>
rect 345 2636 405 2642
rect 345 2614 348 2636
rect 402 2614 405 2636
rect 345 2608 405 2614
rect 425 2639 454 2642
rect 425 2611 431 2639
rect 448 2611 454 2639
rect 382 2581 411 2584
rect 366 2564 388 2581
rect 405 2564 411 2581
rect 382 2561 411 2564
rect 345 2530 405 2536
rect 345 2450 348 2530
rect 402 2450 405 2530
rect 345 2444 405 2450
rect 425 2533 454 2611
rect 425 2447 431 2533
rect 448 2447 454 2533
rect 425 2444 454 2447
<< end >>
