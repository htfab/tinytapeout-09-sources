magic
tech sky130A
magscale 1 2
timestamp 1730822054
<< nwell >>
rect -72 4960 972 5300
rect -72 4908 20 4960
rect 62 4946 108 4960
rect 110 4952 218 4960
rect -72 4296 28 4908
rect -72 4236 20 4296
rect 326 4236 548 4960
rect 854 4236 972 4960
<< pwell >>
rect 226 4120 324 4124
rect -130 2090 1444 4098
<< psubdiff >>
rect -94 3974 2 4060
rect 874 3974 970 4060
rect 874 3378 970 3412
rect 874 3284 986 3378
rect 1294 3284 1408 3378
rect 874 3282 970 3284
rect 2 3202 44 3282
rect 856 3202 970 3282
rect 1312 3254 1408 3284
rect -94 2202 2 2236
rect 1312 2202 1408 2236
rect -94 2090 26 2202
rect 1288 2090 1408 2202
<< nsubdiff >>
rect -34 5106 -10 5264
rect 912 5106 936 5264
rect -34 5072 2 5106
rect -34 4294 2 4318
rect 344 4294 530 4318
rect 872 4294 908 4318
<< psubdiffcont >>
rect 2 4026 874 4060
rect -94 2236 2 3974
rect 416 3282 456 4026
rect 874 3412 970 3974
rect 986 3284 1294 3378
rect 44 3202 856 3282
rect 1312 2236 1408 3254
rect 26 2090 1288 2202
<< nsubdiffcont >>
rect -10 5106 912 5264
rect -34 4318 2 5072
rect 344 4318 530 5106
rect 872 4318 908 5106
<< poly >>
rect 114 5056 206 5072
rect 114 5022 158 5056
rect 192 5022 206 5056
rect 114 5006 206 5022
rect 114 4924 144 5006
rect 668 5056 760 5072
rect 668 5022 682 5056
rect 716 5022 760 5056
rect 668 5006 760 5022
rect 730 4924 760 5006
rect 202 4212 232 4272
rect 642 4260 672 4274
rect 490 4244 672 4260
rect 202 4182 324 4212
rect 490 4210 506 4244
rect 540 4230 672 4244
rect 540 4210 556 4230
rect 490 4194 556 4210
rect 258 4170 324 4182
rect 258 4136 274 4170
rect 308 4136 324 4170
rect 258 4120 324 4136
rect 316 3396 382 3412
rect 316 3362 332 3396
rect 366 3362 382 3396
rect 316 3346 382 3362
rect 114 3316 382 3346
rect 490 3396 556 3412
rect 490 3362 506 3396
rect 540 3362 556 3396
rect 490 3346 556 3362
rect 490 3316 760 3346
rect 1200 3198 1266 3214
rect 1200 3178 1216 3198
rect 818 3164 1216 3178
rect 1250 3164 1266 3198
rect 818 3148 1266 3164
rect 114 2492 144 2496
rect 202 2492 232 2496
rect 114 2476 232 2492
rect 114 2462 156 2476
rect 140 2442 156 2462
rect 190 2462 232 2476
rect 190 2442 206 2462
rect 140 2426 206 2442
rect 290 2378 320 2496
rect 378 2378 408 2496
rect 466 2492 496 2496
rect 554 2492 584 2496
rect 466 2476 584 2492
rect 466 2462 508 2476
rect 492 2442 508 2462
rect 542 2462 584 2476
rect 542 2442 558 2462
rect 492 2426 558 2442
rect 290 2362 408 2378
rect 290 2348 332 2362
rect 316 2328 332 2348
rect 366 2348 408 2362
rect 642 2378 672 2496
rect 730 2378 760 2496
rect 642 2362 760 2378
rect 642 2348 684 2362
rect 366 2328 382 2348
rect 316 2312 382 2328
rect 668 2328 684 2348
rect 718 2348 760 2362
rect 718 2328 734 2348
rect 668 2312 734 2328
<< polycont >>
rect 158 5022 192 5056
rect 682 5022 716 5056
rect 506 4210 540 4244
rect 274 4136 308 4170
rect 332 3362 366 3396
rect 506 3362 540 3396
rect 1216 3164 1250 3198
rect 156 2442 190 2476
rect 508 2442 542 2476
rect 332 2328 366 2362
rect 684 2328 718 2362
<< locali >>
rect -34 5106 -10 5264
rect 912 5106 936 5264
rect -34 5072 2 5106
rect 152 5056 198 5072
rect 152 5022 158 5056
rect 192 5022 198 5056
rect 152 5006 198 5022
rect -34 4294 2 4318
rect 676 5056 722 5072
rect 676 5022 682 5056
rect 716 5022 722 5056
rect 676 5006 722 5022
rect 344 4294 530 4318
rect 872 4294 908 4318
rect 500 4244 546 4260
rect 500 4210 506 4244
rect 540 4210 546 4244
rect 500 4194 546 4210
rect 268 4170 314 4188
rect 268 4136 274 4170
rect 308 4136 314 4170
rect 268 4120 314 4136
rect -94 3974 2 4060
rect 316 3396 382 3402
rect 316 3362 332 3396
rect 366 3362 382 3396
rect 316 3356 382 3362
rect 874 3974 970 4060
rect 490 3396 556 3402
rect 490 3362 506 3396
rect 540 3362 556 3396
rect 490 3356 556 3362
rect 874 3378 970 3412
rect 874 3284 986 3378
rect 1294 3284 1408 3378
rect 874 3282 970 3284
rect 2 3202 44 3282
rect 856 3202 970 3282
rect 1312 3254 1408 3284
rect 1200 3198 1266 3202
rect 1200 3164 1216 3198
rect 1250 3164 1266 3198
rect 1200 3160 1266 3164
rect 140 2476 206 2482
rect 140 2442 156 2476
rect 190 2442 206 2476
rect 140 2436 206 2442
rect 492 2476 558 2482
rect 492 2442 508 2476
rect 542 2442 558 2476
rect 492 2436 558 2442
rect 316 2362 382 2368
rect 316 2328 332 2362
rect 366 2328 382 2362
rect 316 2322 382 2328
rect 668 2362 734 2368
rect 668 2328 684 2362
rect 718 2328 734 2362
rect 668 2322 734 2328
rect -94 2202 2 2236
rect 1312 2202 1408 2236
rect -94 2090 26 2202
rect 1288 2090 1408 2202
<< viali >>
rect -10 5112 912 5258
rect -34 4318 2 5072
rect 158 5022 192 5056
rect 682 5022 716 5056
rect 506 4210 540 4244
rect 274 4136 308 4170
rect -88 2236 -4 3974
rect 332 3362 366 3396
rect 880 3412 964 3974
rect 506 3362 540 3396
rect 1216 3164 1250 3198
rect 156 2442 190 2476
rect 508 2442 542 2476
rect 332 2328 366 2362
rect 684 2328 718 2362
rect 1318 2236 1402 3254
rect 26 2096 1288 2196
<< metal1 >>
rect -514 5410 1768 5446
rect -514 5354 1208 5410
rect 1264 5354 1768 5410
rect -514 5346 1768 5354
rect -514 5258 1768 5264
rect -514 5112 -10 5258
rect 912 5112 1768 5258
rect -514 5106 1768 5112
rect -40 5072 8 5106
rect -206 4854 -142 4860
rect -206 4802 -200 4854
rect -148 4802 -142 4854
rect -206 4796 -142 4802
rect -200 2492 -142 4796
rect -40 4318 -34 5072
rect 2 4318 8 5072
rect 62 4982 108 5106
rect 146 5070 1268 5076
rect 146 5056 1210 5070
rect 146 5022 158 5056
rect 192 5022 682 5056
rect 716 5022 1210 5056
rect 146 5018 1210 5022
rect 1262 5018 1268 5070
rect 146 5016 1268 5018
rect 1204 5012 1268 5016
rect 62 4936 812 4982
rect 62 4898 108 4936
rect 238 4898 284 4936
rect 590 4898 636 4936
rect 766 4898 812 4936
rect -40 4298 8 4318
rect 150 4260 196 4298
rect 150 4254 556 4260
rect 150 4216 496 4254
rect -74 4138 -6 4144
rect -74 4082 -68 4138
rect -12 4082 -6 4138
rect -74 4066 -6 4082
rect 150 4066 196 4216
rect 490 4200 496 4216
rect 550 4200 556 4254
rect 490 4194 556 4200
rect 258 4180 374 4188
rect 258 4126 264 4180
rect 318 4140 374 4180
rect 678 4140 724 4298
rect 318 4126 1112 4140
rect 258 4120 1112 4126
rect 324 4094 1112 4120
rect -74 4020 284 4066
rect -208 2486 -142 2492
rect -208 2432 -202 2486
rect -148 2432 -142 2486
rect -208 2426 -142 2432
rect -94 3974 2 3986
rect -94 2236 -88 3974
rect -4 2236 2 3974
rect 62 3972 108 4020
rect 238 3972 284 4020
rect 324 3396 374 4094
rect 590 3972 636 4094
rect 766 3972 812 4094
rect 874 3974 970 3986
rect 874 3412 880 3974
rect 964 3412 970 3974
rect 1066 3548 1112 4094
rect 1066 3542 1130 3548
rect 1066 3490 1072 3542
rect 1124 3490 1130 3542
rect 1066 3484 1130 3490
rect 150 3308 196 3372
rect 324 3362 332 3396
rect 366 3362 374 3396
rect 324 3350 374 3362
rect 490 3406 556 3412
rect 490 3352 496 3406
rect 550 3352 556 3406
rect 874 3400 970 3412
rect 490 3346 556 3352
rect 150 3262 548 3308
rect 150 3122 196 3262
rect 326 3228 392 3234
rect 326 3174 334 3228
rect 386 3174 392 3228
rect 326 3168 392 3174
rect 326 3122 372 3168
rect 502 3122 548 3262
rect 678 3234 724 3372
rect 658 3228 724 3234
rect 658 3174 666 3228
rect 718 3174 724 3228
rect 658 3168 724 3174
rect 678 3122 724 3168
rect 766 3190 1164 3236
rect 766 3122 812 3190
rect 942 3122 988 3190
rect 1118 3122 1164 3190
rect 1204 3198 1262 5012
rect 1460 4854 1524 4860
rect 1460 4802 1466 4854
rect 1518 4802 1524 4854
rect 1460 4796 1524 4802
rect 1204 3164 1216 3198
rect 1250 3164 1262 3198
rect 1204 3156 1262 3164
rect 1312 3254 1408 3266
rect 62 2284 108 2522
rect 140 2486 206 2492
rect 140 2432 146 2486
rect 200 2432 206 2486
rect 140 2426 206 2432
rect 238 2284 284 2522
rect 316 2372 382 2378
rect 316 2318 322 2372
rect 376 2318 382 2372
rect 316 2312 382 2318
rect 414 2284 460 2522
rect 492 2486 558 2492
rect 492 2432 498 2486
rect 552 2432 558 2486
rect 492 2426 558 2432
rect 590 2284 636 2522
rect 668 2372 734 2378
rect 668 2318 674 2372
rect 728 2318 734 2372
rect 668 2312 734 2318
rect 766 2284 812 2522
rect 62 2238 812 2284
rect -94 2202 2 2236
rect 854 2202 900 2522
rect 1030 2202 1076 2522
rect 1206 2202 1252 2522
rect 1312 2236 1318 3254
rect 1402 2236 1408 3254
rect 1460 2378 1518 4796
rect 1460 2372 1526 2378
rect 1460 2318 1466 2372
rect 1520 2318 1526 2372
rect 1460 2312 1526 2318
rect 1312 2202 1408 2236
rect -514 2196 1768 2202
rect -514 2096 26 2196
rect 1288 2096 1768 2196
rect -514 2090 1768 2096
<< via1 >>
rect 1208 5354 1264 5410
rect -200 4802 -148 4854
rect 1210 5018 1262 5070
rect 496 4244 550 4254
rect -68 4082 -12 4138
rect 496 4210 506 4244
rect 506 4210 540 4244
rect 540 4210 550 4244
rect 496 4200 550 4210
rect 264 4170 318 4180
rect 264 4136 274 4170
rect 274 4136 308 4170
rect 308 4136 318 4170
rect 264 4126 318 4136
rect -202 2432 -148 2486
rect 1072 3490 1124 3542
rect 496 3396 550 3406
rect 496 3362 506 3396
rect 506 3362 540 3396
rect 540 3362 550 3396
rect 496 3352 550 3362
rect 334 3174 386 3228
rect 666 3174 718 3228
rect 1466 4802 1518 4854
rect 146 2476 200 2486
rect 146 2442 156 2476
rect 156 2442 190 2476
rect 190 2442 200 2476
rect 146 2432 200 2442
rect 322 2362 376 2372
rect 322 2328 332 2362
rect 332 2328 366 2362
rect 366 2328 376 2362
rect 322 2318 376 2328
rect 498 2476 552 2486
rect 498 2442 508 2476
rect 508 2442 542 2476
rect 542 2442 552 2476
rect 498 2432 552 2442
rect 674 2362 728 2372
rect 674 2328 684 2362
rect 684 2328 718 2362
rect 718 2328 728 2362
rect 674 2318 728 2328
rect 1466 2318 1520 2372
<< metal2 >>
rect -206 4854 -142 5546
rect 1204 5410 1268 5416
rect 1204 5354 1208 5410
rect 1264 5354 1268 5410
rect 1204 5070 1268 5354
rect 1204 5018 1210 5070
rect 1262 5018 1268 5070
rect 1204 5012 1268 5018
rect -206 4802 -200 4854
rect -148 4802 -142 4854
rect -206 4796 -142 4802
rect 1460 4854 1524 5546
rect 1460 4802 1466 4854
rect 1518 4802 1524 4854
rect 1460 4796 1524 4802
rect 490 4256 556 4260
rect -424 4188 110 4256
rect 490 4254 1738 4256
rect 490 4200 496 4254
rect 550 4200 1738 4254
rect 490 4196 1738 4200
rect -424 2012 -356 4188
rect 42 4180 324 4188
rect -312 4138 -6 4144
rect -312 4082 -68 4138
rect -12 4082 -6 4138
rect 42 4126 264 4180
rect 318 4126 324 4180
rect 42 4120 324 4126
rect -312 4076 -6 4082
rect -312 2012 -244 4076
rect 490 3406 556 4196
rect 1066 3542 1628 3548
rect 1066 3490 1072 3542
rect 1124 3490 1628 3542
rect 1066 3484 1628 3490
rect 490 3352 496 3406
rect 550 3352 556 3406
rect 490 3346 556 3352
rect 326 3228 724 3234
rect 326 3174 334 3228
rect 386 3174 666 3228
rect 718 3174 724 3228
rect 326 3168 724 3174
rect -208 2486 558 2492
rect -208 2432 -202 2486
rect -148 2432 146 2486
rect 200 2432 498 2486
rect 552 2432 558 2486
rect -208 2426 558 2432
rect 316 2372 1526 2378
rect 316 2318 322 2372
rect 376 2318 674 2372
rect 728 2318 1466 2372
rect 1520 2318 1526 2372
rect 316 2312 1526 2318
rect 1562 2012 1628 3484
rect 1672 2012 1738 4196
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_0
timestamp 1730323530
transform 1 0 129 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_1
timestamp 1730323530
transform 1 0 217 0 1 3672
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_2
timestamp 1730323530
transform 1 0 129 0 1 3672
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_3
timestamp 1730323530
transform 1 0 657 0 1 3672
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_4
timestamp 1730323530
transform 1 0 745 0 1 3672
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_5
timestamp 1730323530
transform 1 0 745 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_6
timestamp 1730323530
transform 1 0 217 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_7
timestamp 1730323530
transform 1 0 305 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_8
timestamp 1730323530
transform 1 0 393 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_9
timestamp 1730323530
transform 1 0 1185 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_10
timestamp 1730323530
transform 1 0 569 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_11
timestamp 1730323530
transform 1 0 657 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_12
timestamp 1730323530
transform 1 0 481 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_13
timestamp 1730323530
transform 1 0 833 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_14
timestamp 1730323530
transform 1 0 921 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_15
timestamp 1730323530
transform 1 0 1009 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__nfet_01v8_NM9Y3C  sky130_fd_pr__nfet_01v8_NM9Y3C_16
timestamp 1730323530
transform 1 0 1097 0 1 2822
box -73 -326 73 326
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 745 0 1 4598
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_1
timestamp 1730191042
transform 1 0 129 0 1 4598
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_2
timestamp 1730191042
transform 1 0 217 0 1 4598
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_3
timestamp 1730191042
transform 1 0 657 0 1 4598
box -109 -362 109 362
<< labels >>
rlabel metal2 -206 5482 -142 5546 0 d
port 1 nsew
rlabel metal2 1460 5482 1524 5546 0 nd
port 2 nsew
rlabel metal1 -514 5382 -450 5446 0 clk
port 3 nsew
rlabel metal2 -312 2012 -244 2080 0 out1
port 4 nsew
rlabel metal2 1562 2012 1628 2078 0 out2
port 5 nsew
rlabel metal1 -514 5200 -450 5264 0 VDD
port 6 nsew
rlabel metal1 -514 2138 -450 2202 0 VSS
port 7 nsew
<< end >>
