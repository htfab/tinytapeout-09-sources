magic
tech sky130A
magscale 1 2
timestamp 1730975828
<< locali >>
rect 2254 283 2643 290
rect 2229 256 3934 283
rect 2229 189 2253 256
rect 2229 175 2254 189
rect 2230 -979 2254 175
rect 2615 175 3934 256
rect 2615 137 2664 175
rect 2627 -979 2664 137
rect 2230 -1025 2664 -979
rect 2430 -2216 2906 -2214
rect 2430 -2250 2870 -2216
rect 2904 -2250 2906 -2216
rect 2430 -2251 2906 -2250
rect 2231 -2854 2661 -2815
rect 2231 -3643 2262 -2854
rect 2629 -3621 2661 -2854
rect 2231 -3645 2261 -3643
rect 2233 -3689 2261 -3645
rect 2629 -3689 3937 -3621
rect 2233 -3712 3937 -3689
<< viali >>
rect 2253 189 2615 256
rect 2254 137 2615 189
rect 2254 -979 2627 137
rect 2393 -2251 2430 -2214
rect 2870 -2250 2904 -2216
rect 2262 -3643 2629 -2854
rect 2261 -3689 2629 -3643
<< metal1 >>
rect 2254 283 2627 290
rect 2229 271 2627 283
rect 2229 256 2637 271
rect 3561 269 3650 272
rect 2953 257 3650 269
rect 2229 189 2253 256
rect 2229 175 2254 189
rect 2230 -979 2254 175
rect 2615 160 2637 256
rect 2926 186 3650 257
rect 2615 137 2664 160
rect 2627 -979 2664 137
rect 2778 66 2847 118
rect 2230 -1025 2664 -979
rect 2707 7 2790 13
rect 2926 7 3015 186
rect 3094 66 3163 118
rect 3410 64 3479 116
rect 3265 7 3317 13
rect 3561 9 3650 186
rect 3725 67 3794 119
rect 2707 -51 2790 -45
rect 2233 -1195 2294 -1025
rect 2372 -1135 2441 -1083
rect 2233 -1367 2377 -1195
rect 2237 -1968 2377 -1367
rect 2440 -1927 2611 -1202
rect 2707 -1884 2786 -51
rect 2440 -1961 2623 -1927
rect 2565 -2019 2623 -1961
rect 2707 -1936 2724 -1884
rect 2776 -1936 2786 -1884
rect 2707 -1968 2786 -1936
rect 2840 -1875 3094 7
rect 2840 -1927 2942 -1875
rect 2994 -1927 3094 -1875
rect 2840 -1963 3094 -1927
rect 3159 -45 3265 7
rect 3317 -45 3413 7
rect 3159 -1877 3413 -45
rect 3159 -1929 3257 -1877
rect 3309 -1929 3413 -1877
rect 3159 -1963 3413 -1929
rect 3475 -1868 3729 9
rect 3817 7 3869 13
rect 3475 -1920 3570 -1868
rect 3622 -1920 3729 -1868
rect 3475 -1961 3729 -1920
rect 3788 -45 3817 7
rect 3788 -51 3869 -45
rect 3788 -1898 3867 -51
rect 3788 -1950 3805 -1898
rect 3857 -1950 3867 -1898
rect 3788 -1968 3867 -1950
rect 2307 -2123 2507 -2025
rect 2565 -2084 3795 -2019
rect 2307 -2214 2515 -2123
rect 2307 -2251 2393 -2214
rect 2430 -2251 2515 -2214
rect 2307 -2323 2515 -2251
rect 2307 -2432 2507 -2323
rect 2565 -2479 2623 -2084
rect 3986 -2171 4186 -1971
rect 2864 -2216 2910 -2204
rect 2864 -2250 2870 -2216
rect 2904 -2250 2910 -2216
rect 2864 -2262 2910 -2250
rect 3560 -2206 3636 -2194
rect 3560 -2258 3570 -2206
rect 3622 -2209 3636 -2206
rect 4058 -2209 4103 -2171
rect 3622 -2254 4103 -2209
rect 3622 -2258 3636 -2254
rect 2868 -2377 2905 -2262
rect 3560 -2266 3636 -2258
rect 3978 -2321 4184 -2286
rect 2777 -2437 3797 -2377
rect 3836 -2443 4184 -2321
rect 3794 -2478 3806 -2477
rect 3857 -2478 4184 -2443
rect 2239 -2491 2374 -2485
rect 2239 -2607 2377 -2491
rect 2237 -2654 2377 -2607
rect 2434 -2652 2635 -2479
rect 2711 -2491 2784 -2488
rect 2844 -2489 3093 -2483
rect 2711 -2497 2790 -2491
rect 2711 -2555 2790 -2549
rect 2237 -2808 2288 -2654
rect 2337 -2658 2377 -2654
rect 2368 -2759 2437 -2707
rect 2235 -2815 2288 -2808
rect 2231 -2854 2661 -2815
rect 2231 -3643 2262 -2854
rect 2629 -3621 2661 -2854
rect 2711 -3383 2784 -2555
rect 2711 -3389 2790 -3383
rect 2711 -3447 2790 -3441
rect 2711 -3455 2784 -3447
rect 2844 -3451 3093 -2541
rect 3158 -2484 3407 -2478
rect 3794 -2483 4184 -2478
rect 3158 -3389 3407 -2536
rect 3158 -3441 3256 -3389
rect 3308 -3441 3407 -3389
rect 3158 -3446 3407 -3441
rect 3471 -2493 3720 -2487
rect 3256 -3447 3308 -3446
rect 2777 -3560 2846 -3508
rect 2932 -3613 3004 -3451
rect 3471 -3455 3720 -2545
rect 3867 -2504 4184 -2483
rect 3867 -2535 4044 -2504
rect 3794 -2596 4044 -2535
rect 3794 -3389 3867 -2596
rect 3794 -3441 3811 -3389
rect 3863 -3441 3867 -3389
rect 3794 -3450 3867 -3441
rect 3093 -3559 3162 -3507
rect 3410 -3559 3479 -3507
rect 3557 -3613 3629 -3455
rect 3727 -3559 3796 -3507
rect 2629 -3630 2667 -3621
rect 2231 -3645 2261 -3643
rect 2233 -3689 2261 -3645
rect 2629 -3689 2671 -3630
rect 2233 -3710 2671 -3689
rect 2932 -3685 3629 -3613
rect 2932 -3691 3618 -3685
rect 2233 -3712 2667 -3710
<< via1 >>
rect 2707 -45 2790 7
rect 2724 -1936 2776 -1884
rect 2942 -1927 2994 -1875
rect 3265 -45 3317 7
rect 3257 -1929 3309 -1877
rect 3570 -1920 3622 -1868
rect 3817 -45 3869 7
rect 3805 -1950 3857 -1898
rect 3570 -2258 3622 -2206
rect 2711 -2549 2790 -2497
rect 2844 -2541 3093 -2489
rect 2711 -3441 2790 -3389
rect 3158 -2536 3407 -2484
rect 3256 -3441 3308 -3389
rect 3471 -2545 3720 -2493
rect 3794 -2535 3867 -2483
rect 3811 -3441 3863 -3389
<< metal2 >>
rect 2701 -45 2707 7
rect 2790 1 2796 7
rect 3259 1 3265 7
rect 2790 -39 3265 1
rect 2790 -45 2796 -39
rect 3259 -45 3265 -39
rect 3317 1 3323 7
rect 3811 1 3817 7
rect 3317 -39 3817 1
rect 3317 -45 3323 -39
rect 3811 -45 3817 -39
rect 3869 -45 3875 7
rect 3570 -1868 3622 -1862
rect 2942 -1875 2994 -1869
rect 2724 -1884 2776 -1878
rect 2942 -1933 2994 -1927
rect 3257 -1877 3309 -1871
rect 3570 -1926 3622 -1920
rect 3805 -1898 3857 -1892
rect 2724 -1942 2776 -1936
rect 2729 -2497 2771 -1942
rect 2943 -2489 2993 -1933
rect 3257 -1935 3309 -1929
rect 3257 -2484 3308 -1935
rect 3573 -2194 3618 -1926
rect 3805 -1956 3857 -1950
rect 3560 -2206 3636 -2194
rect 3560 -2258 3570 -2206
rect 3622 -2258 3636 -2206
rect 3560 -2266 3636 -2258
rect 2705 -2549 2711 -2497
rect 2790 -2549 2796 -2497
rect 2838 -2541 2844 -2489
rect 3093 -2541 3099 -2489
rect 3152 -2536 3158 -2484
rect 3407 -2536 3413 -2484
rect 3573 -2493 3618 -2266
rect 3808 -2483 3853 -1956
rect 3465 -2545 3471 -2493
rect 3720 -2545 3726 -2493
rect 3788 -2535 3794 -2483
rect 3867 -2535 3873 -2483
rect 2705 -3441 2711 -3389
rect 2790 -3394 2796 -3389
rect 3250 -3394 3256 -3389
rect 2790 -3436 3256 -3394
rect 2790 -3441 2796 -3436
rect 3250 -3441 3256 -3436
rect 3308 -3394 3314 -3389
rect 3805 -3394 3811 -3389
rect 3308 -3436 3811 -3394
rect 3308 -3441 3314 -3436
rect 3805 -3441 3811 -3436
rect 3863 -3441 3869 -3389
use sky130_fd_pr__nfet_01v8_BBNS5X  XM1
timestamp 1730931944
transform 1 0 3759 0 1 -2970
box -211 -710 211 710
use sky130_fd_pr__pfet_01v8_XGA8MR  XM2
timestamp 1730931944
transform 1 0 3759 0 1 -981
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_648S5X  XM3 ~/Documents/github_project/adc_dac2/mag
timestamp 1730975153
transform 1 0 2406 0 1 -2569
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGASDL  XM4 ~/Documents/github_project/adc_dac2/mag
timestamp 1730931944
transform 1 0 2407 0 1 -1580
box -211 -619 211 619
use sky130_fd_pr__pfet_01v8_XGA8MR  XM5
timestamp 1730931944
transform 1 0 2811 0 1 -981
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM6
timestamp 1730931944
transform 1 0 3127 0 1 -981
box -211 -1219 211 1219
use sky130_fd_pr__pfet_01v8_XGA8MR  XM7
timestamp 1730931944
transform 1 0 3443 0 1 -981
box -211 -1219 211 1219
use sky130_fd_pr__nfet_01v8_BBNS5X  XM8
timestamp 1730931944
transform 1 0 2811 0 1 -2970
box -211 -710 211 710
use sky130_fd_pr__nfet_01v8_BBNS5X  XM9
timestamp 1730931944
transform 1 0 3127 0 1 -2970
box -211 -710 211 710
use sky130_fd_pr__nfet_01v8_BBNS5X  XM10
timestamp 1730931944
transform 1 0 3443 0 1 -2970
box -211 -710 211 710
<< labels >>
flabel metal1 2363 -3387 2563 -3187 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 2282 -7 2482 193 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 2315 -2323 2515 -2123 0 FreeSans 256 0 0 0 ctrl
port 1 nsew
flabel metal1 3986 -2171 4186 -1971 0 FreeSans 256 0 0 0 b
port 3 nsew
flabel metal1 3982 -2500 4182 -2300 0 FreeSans 256 0 0 0 a
port 2 nsew
<< end >>
