magic
tech sky130A
magscale 1 2
timestamp 1730665133
<< locali >>
rect -10130 11328 -9456 11512
rect -7174 11326 -6500 11510
rect -4094 11314 -3420 11498
rect -1092 11322 -418 11506
rect -12670 10156 -12634 10366
rect -12668 7828 -12528 9066
rect -12662 7820 -12534 7828
rect -10356 7814 -9390 7960
rect -7362 7810 -6396 7956
rect -4490 7804 -3524 7950
rect -1422 7812 -456 7958
rect -10108 7510 -9482 7700
rect -7128 7518 -6502 7708
rect -4132 7522 -3506 7712
rect -1102 7526 -476 7716
rect -10396 4010 -9430 4156
rect -7396 4014 -6430 4160
rect -4338 4006 -3372 4152
rect -1342 4004 -376 4150
rect -10122 3712 -9496 3902
rect -7046 3710 -6420 3900
rect -4088 3722 -3462 3912
rect -1136 3710 -510 3900
rect -10400 212 -9434 358
rect -7374 214 -6408 360
rect -4394 214 -3428 360
rect -1378 202 -412 348
<< metal1 >>
rect -12834 11320 -12482 11514
rect -10130 11328 -9456 11512
rect -7174 11326 -6500 11510
rect -12832 10920 -12764 11320
rect -4094 11314 -3420 11498
rect -1092 11322 -418 11506
rect -11112 11222 -10918 11260
rect -11112 11100 -11078 11222
rect -10946 11100 -10918 11222
rect -11112 11074 -10918 11100
rect -8118 11228 -7924 11262
rect -8118 11106 -8092 11228
rect -7960 11106 -7924 11228
rect -8118 11076 -7924 11106
rect -5132 11260 -4926 11266
rect -5132 11074 -5126 11260
rect -4932 11074 -4926 11260
rect -2110 11238 -1916 11260
rect -2110 11116 -2086 11238
rect -1954 11116 -1916 11238
rect -2110 11090 -1916 11116
rect 886 11236 1080 11260
rect 886 11114 916 11236
rect 1048 11114 1080 11236
rect 886 11090 1080 11114
rect -5132 11068 -4926 11074
rect -12836 10592 -12766 10808
rect -12870 10576 -12728 10592
rect -12870 10432 -12858 10576
rect -12742 10432 -12728 10576
rect -12870 10420 -12728 10432
rect -12836 9722 -12766 10420
rect -8812 10220 -8622 10258
rect -8812 10050 -8794 10220
rect -8658 10050 -8622 10220
rect -2836 10232 -2596 10276
rect -8812 10036 -8622 10050
rect -5806 10180 -5616 10204
rect -5806 10010 -5782 10180
rect -5646 10010 -5616 10180
rect -2836 10054 -2798 10232
rect -2642 10054 -2596 10232
rect 190 10258 378 10272
rect 190 10088 216 10258
rect 352 10088 378 10258
rect 190 10056 378 10088
rect -2836 10016 -2596 10054
rect -5806 9982 -5616 10010
rect -12836 9522 -12768 9608
rect -12902 9498 -12712 9522
rect -12902 9328 -12874 9498
rect -12738 9328 -12712 9498
rect -12394 9440 -12254 9824
rect -12902 9300 -12712 9328
rect -12836 8524 -12768 9300
rect -12834 8128 -12766 8410
rect -13052 8122 -12766 8128
rect -13134 8104 -12766 8122
rect -13134 8000 -12976 8104
rect -12840 8000 -12766 8104
rect -13134 7980 -12766 8000
rect -13134 7332 -13002 7980
rect -12668 7828 -12528 9066
rect -10356 7814 -9390 7960
rect -7362 7810 -6396 7956
rect -4490 7804 -3524 7950
rect -1422 7812 -456 7958
rect -12934 7634 -12766 7756
rect -12936 7618 -12764 7634
rect -12936 7514 -12918 7618
rect -12782 7514 -12764 7618
rect -12936 7498 -12764 7514
rect -10108 7510 -9482 7700
rect -7128 7518 -6502 7708
rect -4132 7522 -3506 7712
rect -1102 7526 -476 7716
rect -12934 7388 -12766 7498
rect -12964 7326 -12766 7388
rect -11110 7420 -10916 7452
rect -12964 7208 -12916 7326
rect -11110 7298 -11076 7420
rect -10944 7298 -10916 7420
rect -11110 7270 -10916 7298
rect -13126 7150 -12916 7208
rect -11112 7266 -10916 7270
rect -13126 6792 -12928 7150
rect -11112 7084 -10918 7266
rect -12890 6846 -12764 7062
rect -12890 6826 -12704 6846
rect -12890 6722 -12856 6826
rect -12720 6722 -12704 6826
rect -12890 6710 -12704 6722
rect -12890 6694 -12764 6710
rect -13080 6688 -12764 6694
rect -13126 6634 -12764 6688
rect -13126 6618 -12806 6634
rect -13126 6228 -13028 6618
rect -12962 6398 -12768 6532
rect -12962 6382 -12764 6398
rect -12962 6278 -12916 6382
rect -12780 6278 -12764 6382
rect -12962 6262 -12764 6278
rect -8798 6324 -8648 6340
rect -12962 6176 -12768 6262
rect -12994 6146 -12768 6176
rect -8798 6184 -8782 6324
rect -8670 6184 -8648 6324
rect -2786 6328 -2636 6358
rect -8798 6154 -8648 6184
rect -2786 6188 -2766 6328
rect -2654 6188 -2636 6328
rect -2786 6172 -2636 6188
rect -12994 6012 -12924 6146
rect -13124 5966 -12924 6012
rect -13124 5654 -12930 5966
rect -12886 5764 -12772 5940
rect -12886 5728 -12682 5764
rect -12886 5624 -12842 5728
rect -12706 5624 -12682 5728
rect -12886 5602 -12682 5624
rect -12886 5498 -12772 5602
rect -13044 5484 -12772 5498
rect -13126 5438 -12772 5484
rect -13126 5416 -12850 5438
rect -13126 5080 -12970 5416
rect -12894 5218 -12776 5352
rect -12894 5194 -12698 5218
rect -12894 5090 -12864 5194
rect -12728 5090 -12698 5194
rect -13126 4930 -13008 5080
rect -12894 5056 -12698 5090
rect -12894 5000 -12776 5056
rect -12950 4932 -12776 5000
rect -12950 4854 -12880 4932
rect -13020 4838 -12880 4854
rect -13020 4828 -12906 4838
rect -13042 4808 -12906 4828
rect -13128 4794 -12906 4808
rect -13128 4776 -12990 4794
rect -13128 4388 -13010 4776
rect -12920 4634 -12764 4724
rect -12920 4488 -12880 4634
rect -12790 4488 -12764 4634
rect -12920 4474 -12764 4488
rect -12944 4382 -12764 4474
rect -12944 4292 -12898 4382
rect -12986 4276 -12898 4292
rect -13132 4184 -12898 4276
rect -13132 4134 -12926 4184
rect -13132 3862 -12964 4134
rect -12908 4000 -12766 4094
rect -13132 3752 -13006 3862
rect -12908 3854 -12880 4000
rect -12790 3854 -12766 4000
rect -12670 3994 -12528 5264
rect -10396 4010 -9430 4156
rect -7396 4014 -6430 4160
rect -4338 4006 -3372 4152
rect -1342 4004 -376 4150
rect -12908 3788 -12766 3854
rect -12954 3744 -12766 3788
rect -12954 3654 -12894 3744
rect -10122 3712 -9496 3902
rect -7046 3710 -6420 3900
rect -4088 3722 -3462 3912
rect -1136 3710 -510 3900
rect -12998 3614 -12894 3654
rect -11078 3628 -10930 3638
rect -12998 3612 -12928 3614
rect -13128 3520 -12928 3612
rect -13128 3192 -12964 3520
rect -12836 3472 -12766 3616
rect -11078 3506 -11070 3628
rect -10938 3506 -10930 3628
rect -11078 3500 -10930 3506
rect -8086 3628 -7938 3636
rect -8086 3506 -8078 3628
rect -7946 3506 -7938 3628
rect -8086 3498 -7938 3506
rect -2084 3620 -1930 3634
rect -2084 3498 -2076 3620
rect -1944 3498 -1930 3620
rect -2084 3490 -1930 3498
rect -12912 3396 -12766 3472
rect -12912 3272 -12880 3396
rect -12776 3272 -12766 3396
rect -12912 3194 -12766 3272
rect -12912 3132 -12770 3194
rect -13054 3102 -12770 3132
rect -13054 3092 -12858 3102
rect -13130 3038 -12858 3092
rect -13130 2532 -13028 3038
rect -12930 2796 -12768 2962
rect -12930 2668 -12912 2796
rect -12826 2668 -12768 2796
rect -12930 2594 -12768 2668
rect -12980 2532 -12768 2594
rect -12980 2456 -12918 2532
rect -13026 2420 -12918 2456
rect -13130 2400 -12918 2420
rect -13130 2352 -12958 2400
rect -13130 1994 -12998 2352
rect -12836 2168 -12762 2422
rect -12902 2160 -12762 2168
rect -12916 2140 -12762 2160
rect -12916 2012 -12876 2140
rect -12790 2012 -12762 2140
rect -12916 1988 -12762 2012
rect -12916 1934 -12800 1988
rect -13428 1898 -12800 1934
rect -13432 1884 -12800 1898
rect -13432 1852 -12802 1884
rect -13432 1336 -13354 1852
rect -13132 1766 -13048 1768
rect -13238 1764 -13048 1766
rect -13296 1664 -13048 1764
rect -13296 1524 -13224 1664
rect -13116 1524 -13048 1664
rect -13296 1336 -13048 1524
rect -12928 1680 -12762 1768
rect -12928 1552 -12904 1680
rect -12818 1552 -12762 1680
rect -12928 1384 -12762 1552
rect -12950 1336 -12762 1384
rect -13296 1332 -13064 1336
rect -13296 1224 -13204 1332
rect -12950 1248 -12904 1336
rect -13030 1228 -12904 1248
rect -13426 1184 -13204 1224
rect -13128 1188 -12904 1228
rect -12838 1222 -12756 1224
rect -12670 1222 -12524 1464
rect -13426 800 -13218 1184
rect -13128 1156 -12934 1188
rect -13128 798 -13002 1156
rect -12838 794 -12524 1222
rect -12838 792 -12756 794
rect -12666 760 -12524 794
rect -12670 666 -12524 760
rect -10400 212 -9434 358
rect -7374 214 -6408 360
rect -4394 214 -3428 360
rect -1378 202 -412 348
<< via1 >>
rect -11078 11100 -10946 11222
rect -8092 11106 -7960 11228
rect -5126 11074 -4932 11260
rect -2086 11116 -1954 11238
rect 916 11114 1048 11236
rect -12858 10432 -12742 10576
rect -11774 10432 -11658 10576
rect -8794 10050 -8658 10220
rect -5782 10010 -5646 10180
rect -2798 10054 -2642 10232
rect 216 10088 352 10258
rect -12874 9328 -12738 9498
rect -12976 8000 -12840 8104
rect -12918 7514 -12782 7618
rect -11076 7298 -10944 7420
rect -8098 7296 -7966 7418
rect -5068 7302 -4936 7424
rect -2088 7292 -1934 7436
rect 918 7316 1050 7438
rect -12856 6722 -12720 6826
rect -12916 6278 -12780 6382
rect -11794 6276 -11638 6400
rect -8782 6184 -8670 6324
rect -5762 6190 -5650 6330
rect -2766 6188 -2654 6328
rect 234 6180 346 6320
rect -12842 5624 -12706 5728
rect -12864 5090 -12728 5194
rect -12880 4488 -12790 4634
rect -12880 3854 -12790 4000
rect -11070 3506 -10938 3628
rect -8078 3506 -7946 3628
rect -5094 3492 -4946 3630
rect -2076 3498 -1944 3620
rect 914 3508 1046 3630
rect -12880 3272 -12776 3396
rect -11764 3278 -11660 3402
rect -8768 3048 -8672 3200
rect -5754 2832 -5658 2984
rect -12912 2668 -12826 2796
rect -2768 2598 -2672 2750
rect 256 2292 352 2444
rect -12876 2012 -12790 2140
rect -13224 1524 -13116 1664
rect -12904 1552 -12818 1680
<< metal2 >>
rect -9858 11512 -9614 11530
rect -11106 11414 1114 11512
rect -11108 11314 1114 11414
rect -11108 11260 -10920 11314
rect -11112 11222 -10918 11260
rect -11112 11100 -11078 11222
rect -10946 11100 -10918 11222
rect -11112 11074 -10918 11100
rect -12872 10576 -11644 10594
rect -12872 10432 -12858 10576
rect -12742 10432 -11774 10576
rect -11658 10432 -11644 10576
rect -12872 10418 -11644 10432
rect -12902 9498 -12712 9522
rect -12902 9328 -12874 9498
rect -12738 9328 -12712 9498
rect -12902 9300 -12712 9328
rect -12996 8104 -12824 8120
rect -12996 8000 -12976 8104
rect -12840 8000 -12824 8104
rect -12996 7984 -12824 8000
rect -9858 7836 -9614 11314
rect -8114 11262 -7926 11314
rect -8118 11228 -7924 11262
rect -8118 11106 -8092 11228
rect -7960 11106 -7924 11228
rect -8118 11076 -7924 11106
rect -8812 10220 -8622 10258
rect -8812 10050 -8794 10220
rect -8658 10050 -8622 10220
rect -8812 10036 -8622 10050
rect -6844 7836 -6600 11314
rect -5122 11266 -4934 11314
rect -5132 11260 -4926 11266
rect -5132 11074 -5126 11260
rect -4932 11074 -4926 11260
rect -5132 11068 -4926 11074
rect -5806 10180 -5616 10204
rect -5806 10010 -5782 10180
rect -5646 10010 -5616 10180
rect -5806 9982 -5616 10010
rect -3838 7836 -3594 11314
rect -2104 11260 -1916 11314
rect -2110 11238 -1916 11260
rect -2110 11116 -2086 11238
rect -1954 11116 -1916 11238
rect -2110 11090 -1916 11116
rect -2836 10254 -2596 10276
rect -2836 10030 -2820 10254
rect -2616 10030 -2596 10254
rect -2836 10016 -2596 10030
rect -866 7836 -622 11314
rect 886 11260 1074 11314
rect 886 11236 1080 11260
rect 886 11114 916 11236
rect 1048 11114 1080 11236
rect 886 11090 1080 11114
rect 190 10258 378 10272
rect 190 10088 216 10258
rect 352 10088 378 10258
rect 190 10056 378 10088
rect -11120 7648 1076 7836
rect -12936 7618 -12764 7634
rect -12936 7514 -12918 7618
rect -12782 7514 -12764 7618
rect -11120 7616 1098 7648
rect -12936 7498 -12764 7514
rect -11112 7452 -10940 7616
rect -11112 7420 -10916 7452
rect -11112 7298 -11076 7420
rect -10944 7298 -10916 7420
rect -11112 7268 -10916 7298
rect -11110 7266 -10916 7268
rect -12876 6826 -12704 6846
rect -12876 6722 -12856 6826
rect -12720 6722 -12704 6826
rect -12876 6710 -12704 6722
rect -11810 6400 -11614 6408
rect -12936 6386 -12764 6398
rect -11810 6386 -11794 6400
rect -12936 6382 -11794 6386
rect -12936 6278 -12916 6382
rect -12780 6296 -11794 6382
rect -12780 6278 -12764 6296
rect -12936 6262 -12764 6278
rect -11810 6276 -11794 6296
rect -11638 6276 -11614 6400
rect -11810 6262 -11614 6276
rect -12874 5728 -12682 5764
rect -12874 5624 -12842 5728
rect -12706 5624 -12682 5728
rect -12874 5602 -12682 5624
rect -12890 5208 -12698 5218
rect -12890 5072 -12874 5208
rect -12708 5072 -12698 5208
rect -12890 5056 -12698 5072
rect -12900 4634 -12772 4660
rect -12900 4488 -12880 4634
rect -12790 4488 -12772 4634
rect -12900 4464 -12772 4488
rect -9858 4044 -9614 7616
rect -8102 7436 -7930 7616
rect -8106 7418 -7930 7436
rect -8106 7296 -8098 7418
rect -7966 7296 -7930 7418
rect -8106 7288 -7930 7296
rect -8106 7286 -7952 7288
rect -8798 6324 -8648 6340
rect -8798 6184 -8782 6324
rect -8670 6184 -8648 6324
rect -8798 6154 -8648 6184
rect -6844 4044 -6600 7616
rect -5078 7424 -4906 7616
rect -5078 7302 -5068 7424
rect -4936 7302 -4906 7424
rect -5078 7292 -4906 7302
rect -5078 7290 -4924 7292
rect -5780 6330 -5630 6356
rect -5780 6190 -5762 6330
rect -5650 6190 -5630 6330
rect -5780 6170 -5630 6190
rect -3838 4044 -3594 7616
rect -2096 7436 -1924 7616
rect -2096 7292 -2088 7436
rect -1934 7292 -1924 7436
rect -2096 7288 -1924 7292
rect -2096 7282 -1928 7288
rect -2786 6328 -2636 6358
rect -2786 6188 -2766 6328
rect -2654 6188 -2636 6328
rect -2786 6172 -2636 6188
rect -866 4044 -622 7616
rect 910 7450 1098 7616
rect 908 7438 1098 7450
rect 908 7316 918 7438
rect 1050 7316 1098 7438
rect 908 7314 1098 7316
rect 908 7306 1062 7314
rect 212 6320 362 6338
rect 212 6180 234 6320
rect 346 6180 362 6320
rect 212 6152 362 6180
rect -12898 4000 -12766 4014
rect -12898 3854 -12880 4000
rect -12790 3854 -12766 4000
rect -12898 3828 -12766 3854
rect -11092 3750 1078 4044
rect -11076 3638 -10928 3750
rect -11078 3628 -10928 3638
rect -11078 3506 -11070 3628
rect -10938 3508 -10928 3628
rect -8090 3636 -7942 3750
rect -5096 3636 -4948 3750
rect -8090 3628 -7938 3636
rect -10938 3506 -10930 3508
rect -8090 3506 -8078 3628
rect -7946 3506 -7938 3628
rect -11078 3500 -10930 3506
rect -8086 3498 -7938 3506
rect -5102 3630 -4936 3636
rect -5102 3492 -5094 3630
rect -4946 3492 -4936 3630
rect -2088 3634 -1940 3750
rect 908 3642 1056 3750
rect -2088 3620 -1930 3634
rect -2088 3498 -2076 3620
rect -1944 3498 -1930 3620
rect 904 3630 1058 3642
rect 904 3508 914 3630
rect 1046 3508 1058 3630
rect 904 3498 1058 3508
rect -2088 3492 -1930 3498
rect -5102 3484 -4936 3492
rect -2084 3490 -1930 3492
rect -12894 3396 -12746 3414
rect -12894 3272 -12880 3396
rect -12776 3388 -12746 3396
rect -11782 3402 -11634 3416
rect -11782 3388 -11764 3402
rect -12776 3282 -11764 3388
rect -12776 3272 -12746 3282
rect -12894 3258 -12746 3272
rect -11782 3278 -11764 3282
rect -11660 3278 -11634 3402
rect -11782 3260 -11634 3278
rect -8812 3200 -8656 3216
rect -8812 3048 -8768 3200
rect -8672 3048 -8656 3200
rect -8812 3018 -8656 3048
rect -5782 2984 -5626 3006
rect -5782 2832 -5754 2984
rect -5658 2832 -5626 2984
rect -12930 2796 -12796 2814
rect -5782 2808 -5626 2832
rect -12930 2668 -12912 2796
rect -12826 2668 -12796 2796
rect -12930 2640 -12796 2668
rect -2808 2750 -2652 2770
rect -2808 2598 -2768 2750
rect -2672 2598 -2652 2750
rect -2808 2572 -2652 2598
rect 222 2444 378 2464
rect 222 2292 256 2444
rect 352 2292 378 2444
rect 222 2266 378 2292
rect -12902 2140 -12768 2168
rect -12902 2012 -12876 2140
rect -12790 2012 -12768 2140
rect -12902 1994 -12768 2012
rect -13248 1664 -13068 1686
rect -13248 1524 -13224 1664
rect -13116 1524 -13068 1664
rect -12934 1680 -12800 1710
rect -12934 1552 -12904 1680
rect -12818 1552 -12800 1680
rect -12934 1536 -12800 1552
rect -13248 1506 -13068 1524
<< via2 >>
rect -12874 9328 -12738 9498
rect -12976 8000 -12840 8104
rect -8794 10050 -8658 10220
rect -5782 10010 -5646 10180
rect -2820 10232 -2616 10254
rect -2820 10054 -2798 10232
rect -2798 10054 -2642 10232
rect -2642 10054 -2616 10232
rect -2820 10030 -2616 10054
rect 216 10088 352 10258
rect -12918 7514 -12782 7618
rect -12856 6722 -12720 6826
rect -12842 5624 -12706 5728
rect -12874 5194 -12708 5208
rect -12874 5090 -12864 5194
rect -12864 5090 -12728 5194
rect -12728 5090 -12708 5194
rect -12874 5072 -12708 5090
rect -12880 4488 -12790 4634
rect -8782 6184 -8670 6324
rect -5762 6190 -5650 6330
rect -2766 6188 -2654 6328
rect 234 6180 346 6320
rect -12880 3854 -12790 4000
rect -8768 3048 -8672 3200
rect -5754 2832 -5658 2984
rect -12912 2668 -12826 2796
rect -2768 2598 -2672 2750
rect 256 2292 352 2444
rect -12876 2012 -12790 2140
rect -13224 1524 -13116 1664
rect -12904 1552 -12818 1680
<< metal3 >>
rect -8812 10232 -8622 10258
rect -12864 10220 -8622 10232
rect -12900 10050 -8794 10220
rect -8658 10050 -8622 10220
rect -2836 10254 -2596 10276
rect -12900 10036 -8622 10050
rect -5806 10180 -5616 10204
rect -12900 10032 -8640 10036
rect -12900 9522 -12706 10032
rect -5806 10020 -5782 10180
rect -5832 10010 -5782 10020
rect -5646 10010 -5616 10180
rect -2836 10030 -2820 10254
rect -2616 10030 -2596 10254
rect 190 10258 378 10272
rect 190 10088 216 10258
rect 352 10088 378 10258
rect 190 10056 378 10088
rect -2836 10016 -2596 10030
rect -5832 9982 -5616 10010
rect -12632 9970 -11790 9972
rect -5832 9970 -5618 9982
rect -12632 9964 -5618 9970
rect -12902 9498 -12706 9522
rect -12902 9328 -12874 9498
rect -12738 9328 -12706 9498
rect -12902 9300 -12706 9328
rect -12900 9298 -12706 9300
rect -12634 9778 -5618 9964
rect -12634 9776 -11790 9778
rect -12634 9290 -12406 9776
rect -8902 9742 -5618 9778
rect -2810 9698 -2622 10016
rect -11844 9696 -9020 9698
rect -12282 9646 -9020 9696
rect -5140 9646 -2622 9698
rect -12282 9476 -2622 9646
rect -12634 8124 -12400 9290
rect -12988 8120 -12400 8124
rect -12996 8104 -12400 8120
rect -12996 8000 -12976 8104
rect -12840 8000 -12400 8104
rect -12996 7994 -12400 8000
rect -12996 7984 -12824 7994
rect -12560 7986 -12400 7994
rect -12278 7868 -12194 9476
rect -11844 9452 -2622 9476
rect -2810 9444 -2622 9452
rect 224 9372 362 10056
rect -12066 9368 362 9372
rect -12068 9256 362 9368
rect -12926 7792 -12192 7868
rect -12922 7634 -12780 7792
rect -12936 7618 -12764 7634
rect -12936 7514 -12918 7618
rect -12782 7514 -12764 7618
rect -12936 7498 -12764 7514
rect -12876 6826 -12704 6846
rect -12876 6722 -12856 6826
rect -12720 6824 -12704 6826
rect -12068 6824 -11962 9256
rect -12720 6722 -11962 6824
rect -12876 6718 -11962 6722
rect -12876 6710 -12704 6718
rect -12068 6714 -11962 6718
rect -8798 6324 -8648 6340
rect -8798 6210 -8782 6324
rect -12720 6184 -8782 6210
rect -8670 6184 -8648 6324
rect -12720 6154 -8648 6184
rect -5780 6330 -5630 6356
rect -5780 6190 -5762 6330
rect -5650 6190 -5630 6330
rect -5780 6170 -5630 6190
rect -2786 6328 -2636 6358
rect -2786 6188 -2766 6328
rect -2654 6188 -2636 6328
rect -2786 6172 -2636 6188
rect 212 6320 362 6338
rect 212 6180 234 6320
rect 346 6180 362 6320
rect -12720 6128 -8666 6154
rect -12716 5764 -12634 6128
rect -8772 6126 -8668 6128
rect -5776 6040 -5632 6170
rect -12874 5758 -12634 5764
rect -12564 5936 -5630 6040
rect -12874 5728 -12632 5758
rect -12874 5624 -12842 5728
rect -12706 5624 -12632 5728
rect -12874 5610 -12632 5624
rect -12874 5606 -12634 5610
rect -12874 5602 -12682 5606
rect -12890 5210 -12698 5218
rect -12564 5210 -12438 5936
rect -2764 5826 -2650 6172
rect 212 6152 362 6180
rect -12314 5822 -2636 5826
rect -12318 5704 -2636 5822
rect -12890 5208 -12432 5210
rect -12890 5072 -12874 5208
rect -12708 5100 -12432 5208
rect -12708 5072 -12698 5100
rect -12564 5098 -12438 5100
rect -12890 5056 -12698 5072
rect -12900 4648 -12772 4660
rect -12318 4648 -12204 5704
rect 248 5600 334 6152
rect -12900 4634 -12204 4648
rect -12900 4488 -12880 4634
rect -12790 4526 -12204 4634
rect -12112 5524 334 5600
rect -12112 5502 330 5524
rect -12790 4488 -12772 4526
rect -12900 4464 -12772 4488
rect -12898 4008 -12766 4014
rect -12112 4008 -12008 5502
rect -12898 4000 -12008 4008
rect -12898 3854 -12880 4000
rect -12790 3916 -12008 4000
rect -12790 3914 -12010 3916
rect -12790 3854 -12766 3914
rect -12898 3828 -12766 3854
rect -8812 3200 -8656 3216
rect -8812 3184 -8768 3200
rect -12922 3172 -8768 3184
rect -12926 3084 -8768 3172
rect -12926 2814 -12822 3084
rect -8812 3048 -8768 3084
rect -8672 3048 -8656 3200
rect -8812 3018 -8656 3048
rect -5782 2984 -5626 3006
rect -5782 2936 -5754 2984
rect -12706 2920 -5754 2936
rect -12710 2832 -5754 2920
rect -5658 2832 -5626 2984
rect -12930 2796 -12796 2814
rect -12710 2808 -5626 2832
rect -12710 2804 -5642 2808
rect -12930 2668 -12912 2796
rect -12826 2668 -12796 2796
rect -12930 2640 -12796 2668
rect -12902 2140 -12768 2168
rect -12902 2012 -12876 2140
rect -12790 2130 -12768 2140
rect -12706 2130 -12598 2804
rect -2808 2750 -2652 2770
rect -2808 2706 -2768 2750
rect -12464 2598 -2768 2706
rect -2672 2598 -2652 2750
rect -12464 2576 -2652 2598
rect -12790 2016 -12598 2130
rect -12790 2012 -12768 2016
rect -12902 1994 -12768 2012
rect -12706 2010 -12598 2016
rect -12460 1886 -12330 2576
rect -2808 2572 -2652 2576
rect 222 2444 378 2464
rect 222 2408 256 2444
rect -13238 1774 -12330 1886
rect -12224 2312 256 2408
rect -13234 1686 -13112 1774
rect -12934 1694 -12800 1710
rect -12224 1694 -12114 2312
rect 222 2292 256 2312
rect 352 2292 378 2444
rect 222 2266 378 2292
rect -13248 1664 -13068 1686
rect -13248 1524 -13224 1664
rect -13116 1524 -13068 1664
rect -12934 1680 -12114 1694
rect -12934 1552 -12904 1680
rect -12818 1556 -12114 1680
rect -12818 1552 -12800 1556
rect -12934 1536 -12800 1552
rect -12224 1538 -12114 1556
rect -13248 1506 -13068 1524
use compr0  compr0_0
timestamp 1730635755
transform 1 0 -1832 0 1 596
box 1230 -398 4034 3312
use compr1  compr1_0
timestamp 1730635755
transform 1 0 -1828 0 1 4402
box 1230 -398 4034 3312
use compr2  compr2_0
timestamp 1730635755
transform 1 0 -1832 0 1 8196
box 1230 -398 4034 3312
use compr3  compr3_0
timestamp 1730635755
transform 1 0 -4824 0 1 596
box 1230 -398 4034 3312
use compr4  compr4_0
timestamp 1730635755
transform 1 0 -4830 0 1 4396
box 1230 -398 4034 3312
use compr5  compr5_0
timestamp 1730635755
transform 1 0 -4830 0 1 8196
box 1230 -398 4034 3312
use compr6  compr6_0
timestamp 1730635755
transform 1 0 -7832 0 1 596
box 1230 -398 4034 3312
use compr7  compr7_0
timestamp 1730635755
transform 1 0 -7826 0 1 4396
box 1230 -398 4034 3312
use compr8  compr8_0
timestamp 1730635755
transform 1 0 -7832 0 1 8196
box 1230 -398 4034 3312
use compr9  compr9_0
timestamp 1730635755
transform 1 0 -10834 0 1 596
box 1230 -398 4034 3312
use compr10  compr10_0
timestamp 1730635755
transform 1 0 -10834 0 1 4396
box 1230 -398 4034 3312
use compr11  compr11_0
timestamp 1730635755
transform 1 0 -10834 0 1 8196
box 1230 -398 4034 3312
use compr12  compr12_0
timestamp 1730635755
transform 1 0 -13822 0 1 596
box 1230 -398 4034 3312
use compr13  compr13_0
timestamp 1730635755
transform 1 0 -13830 0 1 4398
box 1230 -398 4034 3312
use compr14  compr14_0
timestamp 1730635755
transform 1 0 -13830 0 1 8200
box 1230 -398 4034 3312
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR1
timestamp 1730493024
transform 1 0 -12801 0 1 1280
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730493024
transform 1 0 -12801 0 1 7270
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR3
timestamp 1730493024
transform 1 0 -12801 0 1 10864
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR4
timestamp 1730493024
transform 1 0 -13393 0 1 1280
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR5
timestamp 1730493024
transform 1 0 -12801 0 1 8468
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730493024
transform 1 0 -13097 0 1 7270
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR7
timestamp 1730493024
transform 1 0 -12801 0 1 9666
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730493024
transform 1 0 -13097 0 1 4874
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR9
timestamp 1730493024
transform 1 0 -12801 0 1 2478
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730493024
transform 1 0 -13097 0 1 3676
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR11
timestamp 1730493024
transform 1 0 -13097 0 1 1280
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730493024
transform 1 0 -13097 0 1 2478
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR13
timestamp 1730493024
transform 1 0 -12801 0 1 3676
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730493024
transform 1 0 -12801 0 1 4874
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR15
timestamp 1730493024
transform 1 0 -12801 0 1 6072
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730493024
transform 1 0 -13097 0 1 6072
box -201 -652 201 652
<< end >>
