magic
tech sky130A
magscale 1 2
timestamp 1730975153
<< error_p >>
rect -29 431 29 437
rect -29 397 -17 431
rect -29 391 29 397
rect -29 -397 29 -391
rect -29 -431 -17 -397
rect -29 -437 29 -431
<< nwell >>
rect -211 -569 211 569
<< pmos >>
rect -15 -350 15 350
<< pdiff >>
rect -73 338 -15 350
rect -73 -338 -61 338
rect -27 -338 -15 338
rect -73 -350 -15 -338
rect 15 338 73 350
rect 15 -338 27 338
rect 61 -338 73 338
rect 15 -350 73 -338
<< pdiffc >>
rect -61 -338 -27 338
rect 27 -338 61 338
<< nsubdiff >>
rect -175 499 -79 533
rect 79 499 175 533
rect -175 437 -141 499
rect 141 437 175 499
rect -175 -499 -141 -437
rect 141 -499 175 -437
rect -175 -533 -79 -499
rect 79 -533 175 -499
<< nsubdiffcont >>
rect -79 499 79 533
rect -175 -437 -141 437
rect 141 -437 175 437
rect -79 -533 79 -499
<< poly >>
rect -33 431 33 447
rect -33 397 -17 431
rect 17 397 33 431
rect -33 381 33 397
rect -15 350 15 381
rect -15 -381 15 -350
rect -33 -397 33 -381
rect -33 -431 -17 -397
rect 17 -431 33 -397
rect -33 -447 33 -431
<< polycont >>
rect -17 397 17 431
rect -17 -431 17 -397
<< locali >>
rect -175 499 -79 533
rect 79 499 175 533
rect -175 437 -141 499
rect 141 437 175 499
rect -33 397 -17 431
rect 17 397 33 431
rect -61 338 -27 354
rect -61 -354 -27 -338
rect 27 338 61 354
rect 27 -354 61 -338
rect -33 -431 -17 -397
rect 17 -431 33 -397
rect -175 -499 -141 -437
rect 141 -499 175 -437
rect -175 -533 -79 -499
rect 79 -533 175 -499
<< viali >>
rect -17 397 17 431
rect -61 -338 -27 338
rect 27 -338 61 338
rect -17 -431 17 -397
<< metal1 >>
rect -29 431 29 437
rect -29 397 -17 431
rect 17 397 29 431
rect -29 391 29 397
rect -67 338 -21 350
rect -67 -338 -61 338
rect -27 -338 -21 338
rect -67 -350 -21 -338
rect 21 338 67 350
rect 21 -338 27 338
rect 61 -338 67 338
rect 21 -350 67 -338
rect -29 -397 29 -391
rect -29 -431 -17 -397
rect 17 -431 29 -397
rect -29 -437 29 -431
<< properties >>
string FIXED_BBOX -158 -516 158 516
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
