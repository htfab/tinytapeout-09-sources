magic
tech sky130A
magscale 1 2
timestamp 1730749971
<< nwell >>
rect 30 954 428 1086
rect 30 230 120 954
rect 338 896 428 954
rect 328 288 428 896
rect 338 230 428 288
<< pwell >>
rect 30 -196 428 230
<< psubdiff >>
rect 66 142 102 166
rect 66 -100 102 -64
rect 356 142 392 166
rect 356 -100 392 -64
rect 66 -196 104 -100
rect 354 -196 392 -100
<< nsubdiff >>
rect 66 954 104 1050
rect 354 954 392 1050
rect 66 920 102 954
rect 66 288 102 312
rect 356 920 392 954
rect 356 288 392 312
<< psubdiffcont >>
rect 66 -64 102 142
rect 356 -64 392 142
rect 104 -196 354 -100
<< nsubdiffcont >>
rect 104 954 354 1050
rect 66 312 102 920
rect 356 312 392 920
<< poly >>
rect 214 254 244 266
rect 136 244 244 254
rect 136 210 152 244
rect 190 210 244 244
rect 136 200 244 210
rect 214 188 244 200
<< polycont >>
rect 152 210 190 244
<< locali >>
rect 66 954 104 1050
rect 354 954 392 1050
rect 66 920 102 954
rect 66 288 102 312
rect 356 920 392 954
rect 356 288 392 312
rect 136 244 206 254
rect 136 210 152 244
rect 190 210 206 244
rect 136 200 206 210
rect 66 142 102 166
rect 66 -100 102 -64
rect 356 142 392 166
rect 356 -100 392 -64
rect 66 -196 104 -100
rect 354 -196 392 -100
<< viali >>
rect 104 962 354 1042
rect 66 312 102 920
rect 356 312 392 920
rect 152 210 190 244
rect 66 -64 102 142
rect 356 -64 392 142
rect 104 -188 354 -108
<< metal1 >>
rect 30 1042 428 1050
rect 30 962 104 1042
rect 354 962 428 1042
rect 30 954 428 962
rect 60 920 108 954
rect 60 312 66 920
rect 102 312 108 920
rect 162 892 208 954
rect 350 920 398 954
rect 60 288 108 312
rect 350 312 356 920
rect 392 312 398 920
rect 136 244 206 254
rect 136 210 152 244
rect 190 210 206 244
rect 136 200 206 210
rect 60 142 108 166
rect 250 162 296 292
rect 350 288 398 312
rect 60 -64 66 142
rect 102 -64 108 142
rect 350 142 398 166
rect 60 -100 108 -64
rect 162 -100 208 -38
rect 350 -64 356 142
rect 392 -64 398 142
rect 350 -100 398 -64
rect 30 -108 428 -100
rect 30 -188 104 -108
rect 354 -188 428 -108
rect 30 -196 428 -188
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1730191042
transform 1 0 229 0 1 62
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 229 0 1 592
box -109 -362 109 362
<< end >>
