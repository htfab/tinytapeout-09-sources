** sch_path: /home/ttuser/Desktop/tt09-sar-adc-dac-combo/xschem/dacswitch.sch
.subckt dacswitch GND VDDA Cin VDD VOUT
*.PININFO GND:B VDDA:B Cin:I VDD:B VOUT:O
x3 net5 VGND VNB VPB VPWR net4 sky130_fd_sc_hd__inv_1
x4 Cin net3 VGND VNB VPB VPWR VOUT sky130_fd_sc_hd__nor2_1
x5 Cin VGND VNB VPB VPWR net1 sky130_fd_sc_hd__inv_1
x6 net4 net1 VGND VNB VPB VPWR net2 sky130_fd_sc_hd__nor2_1
x7 VOUT VGND VNB VPB VPWR net5 sky130_fd_sc_hd__inv_1
x8 net6 VGND VNB VPB VPWR net3 sky130_fd_sc_hd__inv_1
x9 net2 VGND VNB VPB VPWR net6 sky130_fd_sc_hd__inv_1
.ends
.end
