magic
tech sky130A
magscale 1 2
timestamp 1728214159
<< error_p >>
rect -365 2081 -307 2087
rect -173 2081 -115 2087
rect 19 2081 77 2087
rect 211 2081 269 2087
rect 403 2081 461 2087
rect -365 2047 -353 2081
rect -173 2047 -161 2081
rect 19 2047 31 2081
rect 211 2047 223 2081
rect 403 2047 415 2081
rect -365 2041 -307 2047
rect -173 2041 -115 2047
rect 19 2041 77 2047
rect 211 2041 269 2047
rect 403 2041 461 2047
rect -461 -2047 -403 -2041
rect -269 -2047 -211 -2041
rect -77 -2047 -19 -2041
rect 115 -2047 173 -2041
rect 307 -2047 365 -2041
rect -461 -2081 -449 -2047
rect -269 -2081 -257 -2047
rect -77 -2081 -65 -2047
rect 115 -2081 127 -2047
rect 307 -2081 319 -2047
rect -461 -2087 -403 -2081
rect -269 -2087 -211 -2081
rect -77 -2087 -19 -2081
rect 115 -2087 173 -2081
rect 307 -2087 365 -2081
<< nwell >>
rect -647 -2219 647 2219
<< pmos >>
rect -447 -2000 -417 2000
rect -351 -2000 -321 2000
rect -255 -2000 -225 2000
rect -159 -2000 -129 2000
rect -63 -2000 -33 2000
rect 33 -2000 63 2000
rect 129 -2000 159 2000
rect 225 -2000 255 2000
rect 321 -2000 351 2000
rect 417 -2000 447 2000
<< pdiff >>
rect -509 1988 -447 2000
rect -509 -1988 -497 1988
rect -463 -1988 -447 1988
rect -509 -2000 -447 -1988
rect -417 1988 -351 2000
rect -417 -1988 -401 1988
rect -367 -1988 -351 1988
rect -417 -2000 -351 -1988
rect -321 1988 -255 2000
rect -321 -1988 -305 1988
rect -271 -1988 -255 1988
rect -321 -2000 -255 -1988
rect -225 1988 -159 2000
rect -225 -1988 -209 1988
rect -175 -1988 -159 1988
rect -225 -2000 -159 -1988
rect -129 1988 -63 2000
rect -129 -1988 -113 1988
rect -79 -1988 -63 1988
rect -129 -2000 -63 -1988
rect -33 1988 33 2000
rect -33 -1988 -17 1988
rect 17 -1988 33 1988
rect -33 -2000 33 -1988
rect 63 1988 129 2000
rect 63 -1988 79 1988
rect 113 -1988 129 1988
rect 63 -2000 129 -1988
rect 159 1988 225 2000
rect 159 -1988 175 1988
rect 209 -1988 225 1988
rect 159 -2000 225 -1988
rect 255 1988 321 2000
rect 255 -1988 271 1988
rect 305 -1988 321 1988
rect 255 -2000 321 -1988
rect 351 1988 417 2000
rect 351 -1988 367 1988
rect 401 -1988 417 1988
rect 351 -2000 417 -1988
rect 447 1988 509 2000
rect 447 -1988 463 1988
rect 497 -1988 509 1988
rect 447 -2000 509 -1988
<< pdiffc >>
rect -497 -1988 -463 1988
rect -401 -1988 -367 1988
rect -305 -1988 -271 1988
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
rect 271 -1988 305 1988
rect 367 -1988 401 1988
rect 463 -1988 497 1988
<< nsubdiff >>
rect -611 2149 -515 2183
rect 515 2149 611 2183
rect -611 2087 -577 2149
rect 577 2087 611 2149
rect -611 -2149 -577 -2087
rect 577 -2149 611 -2087
rect -611 -2183 -515 -2149
rect 515 -2183 611 -2149
<< nsubdiffcont >>
rect -515 2149 515 2183
rect -611 -2087 -577 2087
rect 577 -2087 611 2087
rect -515 -2183 515 -2149
<< poly >>
rect -369 2081 -303 2097
rect -369 2047 -353 2081
rect -319 2047 -303 2081
rect -369 2031 -303 2047
rect -177 2081 -111 2097
rect -177 2047 -161 2081
rect -127 2047 -111 2081
rect -177 2031 -111 2047
rect 15 2081 81 2097
rect 15 2047 31 2081
rect 65 2047 81 2081
rect 15 2031 81 2047
rect 207 2081 273 2097
rect 207 2047 223 2081
rect 257 2047 273 2081
rect 207 2031 273 2047
rect 399 2081 465 2097
rect 399 2047 415 2081
rect 449 2047 465 2081
rect 399 2031 465 2047
rect -447 2000 -417 2026
rect -351 2000 -321 2031
rect -255 2000 -225 2026
rect -159 2000 -129 2031
rect -63 2000 -33 2026
rect 33 2000 63 2031
rect 129 2000 159 2026
rect 225 2000 255 2031
rect 321 2000 351 2026
rect 417 2000 447 2031
rect -447 -2031 -417 -2000
rect -351 -2026 -321 -2000
rect -255 -2031 -225 -2000
rect -159 -2026 -129 -2000
rect -63 -2031 -33 -2000
rect 33 -2026 63 -2000
rect 129 -2031 159 -2000
rect 225 -2026 255 -2000
rect 321 -2031 351 -2000
rect 417 -2026 447 -2000
rect -465 -2047 -399 -2031
rect -465 -2081 -449 -2047
rect -415 -2081 -399 -2047
rect -465 -2097 -399 -2081
rect -273 -2047 -207 -2031
rect -273 -2081 -257 -2047
rect -223 -2081 -207 -2047
rect -273 -2097 -207 -2081
rect -81 -2047 -15 -2031
rect -81 -2081 -65 -2047
rect -31 -2081 -15 -2047
rect -81 -2097 -15 -2081
rect 111 -2047 177 -2031
rect 111 -2081 127 -2047
rect 161 -2081 177 -2047
rect 111 -2097 177 -2081
rect 303 -2047 369 -2031
rect 303 -2081 319 -2047
rect 353 -2081 369 -2047
rect 303 -2097 369 -2081
<< polycont >>
rect -353 2047 -319 2081
rect -161 2047 -127 2081
rect 31 2047 65 2081
rect 223 2047 257 2081
rect 415 2047 449 2081
rect -449 -2081 -415 -2047
rect -257 -2081 -223 -2047
rect -65 -2081 -31 -2047
rect 127 -2081 161 -2047
rect 319 -2081 353 -2047
<< locali >>
rect -611 2149 -515 2183
rect 515 2149 611 2183
rect -611 2087 -577 2149
rect 577 2087 611 2149
rect -369 2047 -353 2081
rect -319 2047 -303 2081
rect -177 2047 -161 2081
rect -127 2047 -111 2081
rect 15 2047 31 2081
rect 65 2047 81 2081
rect 207 2047 223 2081
rect 257 2047 273 2081
rect 399 2047 415 2081
rect 449 2047 465 2081
rect -497 1988 -463 2004
rect -497 -2004 -463 -1988
rect -401 1988 -367 2004
rect -401 -2004 -367 -1988
rect -305 1988 -271 2004
rect -305 -2004 -271 -1988
rect -209 1988 -175 2004
rect -209 -2004 -175 -1988
rect -113 1988 -79 2004
rect -113 -2004 -79 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 79 1988 113 2004
rect 79 -2004 113 -1988
rect 175 1988 209 2004
rect 175 -2004 209 -1988
rect 271 1988 305 2004
rect 271 -2004 305 -1988
rect 367 1988 401 2004
rect 367 -2004 401 -1988
rect 463 1988 497 2004
rect 463 -2004 497 -1988
rect -465 -2081 -449 -2047
rect -415 -2081 -399 -2047
rect -273 -2081 -257 -2047
rect -223 -2081 -207 -2047
rect -81 -2081 -65 -2047
rect -31 -2081 -15 -2047
rect 111 -2081 127 -2047
rect 161 -2081 177 -2047
rect 303 -2081 319 -2047
rect 353 -2081 369 -2047
rect -611 -2149 -577 -2087
rect 577 -2149 611 -2087
rect -611 -2183 -515 -2149
rect 515 -2183 611 -2149
<< viali >>
rect -353 2047 -319 2081
rect -161 2047 -127 2081
rect 31 2047 65 2081
rect 223 2047 257 2081
rect 415 2047 449 2081
rect -497 -1988 -463 1988
rect -401 -1988 -367 1988
rect -305 -1988 -271 1988
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
rect 271 -1988 305 1988
rect 367 -1988 401 1988
rect 463 -1988 497 1988
rect -449 -2081 -415 -2047
rect -257 -2081 -223 -2047
rect -65 -2081 -31 -2047
rect 127 -2081 161 -2047
rect 319 -2081 353 -2047
<< metal1 >>
rect -365 2081 -307 2087
rect -365 2047 -353 2081
rect -319 2047 -307 2081
rect -365 2041 -307 2047
rect -173 2081 -115 2087
rect -173 2047 -161 2081
rect -127 2047 -115 2081
rect -173 2041 -115 2047
rect 19 2081 77 2087
rect 19 2047 31 2081
rect 65 2047 77 2081
rect 19 2041 77 2047
rect 211 2081 269 2087
rect 211 2047 223 2081
rect 257 2047 269 2081
rect 211 2041 269 2047
rect 403 2081 461 2087
rect 403 2047 415 2081
rect 449 2047 461 2081
rect 403 2041 461 2047
rect -503 1988 -457 2000
rect -503 -1988 -497 1988
rect -463 -1988 -457 1988
rect -503 -2000 -457 -1988
rect -407 1988 -361 2000
rect -407 -1988 -401 1988
rect -367 -1988 -361 1988
rect -407 -2000 -361 -1988
rect -311 1988 -265 2000
rect -311 -1988 -305 1988
rect -271 -1988 -265 1988
rect -311 -2000 -265 -1988
rect -215 1988 -169 2000
rect -215 -1988 -209 1988
rect -175 -1988 -169 1988
rect -215 -2000 -169 -1988
rect -119 1988 -73 2000
rect -119 -1988 -113 1988
rect -79 -1988 -73 1988
rect -119 -2000 -73 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 73 1988 119 2000
rect 73 -1988 79 1988
rect 113 -1988 119 1988
rect 73 -2000 119 -1988
rect 169 1988 215 2000
rect 169 -1988 175 1988
rect 209 -1988 215 1988
rect 169 -2000 215 -1988
rect 265 1988 311 2000
rect 265 -1988 271 1988
rect 305 -1988 311 1988
rect 265 -2000 311 -1988
rect 361 1988 407 2000
rect 361 -1988 367 1988
rect 401 -1988 407 1988
rect 361 -2000 407 -1988
rect 457 1988 503 2000
rect 457 -1988 463 1988
rect 497 -1988 503 1988
rect 457 -2000 503 -1988
rect -461 -2047 -403 -2041
rect -461 -2081 -449 -2047
rect -415 -2081 -403 -2047
rect -461 -2087 -403 -2081
rect -269 -2047 -211 -2041
rect -269 -2081 -257 -2047
rect -223 -2081 -211 -2047
rect -269 -2087 -211 -2081
rect -77 -2047 -19 -2041
rect -77 -2081 -65 -2047
rect -31 -2081 -19 -2047
rect -77 -2087 -19 -2081
rect 115 -2047 173 -2041
rect 115 -2081 127 -2047
rect 161 -2081 173 -2047
rect 115 -2087 173 -2081
rect 307 -2047 365 -2041
rect 307 -2081 319 -2047
rect 353 -2081 365 -2047
rect 307 -2087 365 -2081
<< properties >>
string FIXED_BBOX -594 -2166 594 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
