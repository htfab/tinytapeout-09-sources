** sch_path: /home/ttuser/Desktop/tt09-sar-adc-dac-combo/xschem/lthinverter.sch
.subckt lthinverter VDDA GND VOUT VIN
*.PININFO VOUT:O GND:B VIN:I VDDA:B
XM9 VOUT VIN VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM3 VOUT VIN GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends
.GLOBAL GND
.GLOBAL VDDA
.end
