magic
tech sky130A
magscale 1 2
timestamp 1730892491
<< error_p >>
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
<< nwell >>
rect -211 -719 211 719
<< pmos >>
rect -15 -500 15 500
<< pdiff >>
rect -73 488 -15 500
rect -73 -488 -61 488
rect -27 -488 -15 488
rect -73 -500 -15 -488
rect 15 488 73 500
rect 15 -488 27 488
rect 61 -488 73 488
rect 15 -500 73 -488
<< pdiffc >>
rect -61 -488 -27 488
rect 27 -488 61 488
<< nsubdiff >>
rect -175 649 -79 683
rect 79 649 175 683
rect -175 587 -141 649
rect 141 587 175 649
rect -175 -649 -141 -587
rect 141 -649 175 -587
rect -175 -683 -79 -649
rect 79 -683 175 -649
<< nsubdiffcont >>
rect -79 649 79 683
rect -175 -587 -141 587
rect 141 -587 175 587
rect -79 -683 79 -649
<< poly >>
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -15 500 15 531
rect -15 -531 15 -500
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
<< polycont >>
rect -17 547 17 581
rect -17 -581 17 -547
<< locali >>
rect -175 649 -79 683
rect 79 649 175 683
rect -175 587 -141 649
rect 141 587 175 649
rect -33 547 -17 581
rect 17 547 33 581
rect -61 488 -27 504
rect -61 -504 -27 -488
rect 27 488 61 504
rect 27 -504 61 -488
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -175 -649 -141 -587
rect 141 -649 175 -587
rect -175 -683 -79 -649
rect 79 -683 175 -649
<< viali >>
rect -17 547 17 581
rect -61 -488 -27 488
rect 27 -488 61 488
rect -17 -581 17 -547
<< metal1 >>
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -67 488 -21 500
rect -67 -488 -61 488
rect -27 -488 -21 488
rect -67 -500 -21 -488
rect 21 488 67 500
rect 21 -488 27 488
rect 61 -488 67 488
rect 21 -500 67 -488
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
<< properties >>
string FIXED_BBOX -158 -666 158 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
