magic
tech sky130A
magscale 1 2
timestamp 1731228565
<< nwell >>
rect 348 860 1260 1814
<< pwell >>
rect 348 -416 1260 860
<< psubdiff >>
rect 450 794 516 834
rect 1156 794 1228 834
rect 450 758 490 794
rect 1188 764 1228 794
rect 450 130 490 164
rect 450 90 516 130
rect 658 90 720 130
rect 680 60 720 90
rect 680 -272 720 -238
rect 1188 -272 1228 -238
rect 388 -416 412 -272
rect 1228 -416 1252 -272
<< nsubdiff >>
rect 384 1634 414 1778
rect 1200 1634 1224 1778
rect 538 1600 578 1634
rect 538 976 578 1000
rect 832 1600 930 1634
rect 832 976 930 1000
rect 1184 1600 1224 1634
rect 1184 974 1224 1000
<< psubdiffcont >>
rect 516 794 1156 834
rect 450 164 490 758
rect 516 90 658 130
rect 680 -238 720 60
rect 1188 -238 1228 764
rect 412 -416 1228 -272
<< nsubdiffcont >>
rect 414 1634 1200 1778
rect 538 1000 578 1600
rect 832 1000 930 1600
rect 1184 1000 1224 1600
<< poly >>
rect 690 938 720 954
rect 626 928 720 938
rect 1042 936 1072 952
rect 626 894 642 928
rect 676 894 720 928
rect 626 884 720 894
rect 978 926 1072 936
rect 978 892 994 926
rect 1028 892 1072 926
rect 978 882 1072 892
rect 978 746 1072 756
rect 978 712 994 746
rect 1028 712 1072 746
rect 978 702 1072 712
rect 1042 660 1072 702
rect 602 378 984 408
rect 722 368 776 378
rect 722 334 732 368
rect 766 334 776 368
rect 722 318 776 334
rect 954 326 1140 336
rect 954 306 1090 326
rect 1074 292 1090 306
rect 1124 292 1140 326
rect 1074 282 1140 292
rect 866 -158 896 -146
rect 854 -174 908 -158
rect 854 -208 864 -174
rect 898 -208 908 -174
rect 854 -224 908 -208
<< polycont >>
rect 642 894 676 928
rect 994 892 1028 926
rect 994 712 1028 746
rect 732 334 766 368
rect 1090 292 1124 326
rect 864 -208 898 -174
<< locali >>
rect 384 1634 414 1778
rect 1200 1634 1224 1778
rect 538 1600 578 1634
rect 538 976 578 1000
rect 832 1600 930 1634
rect 832 976 930 1000
rect 1184 1600 1224 1634
rect 1184 974 1224 1000
rect 626 928 692 938
rect 626 894 642 928
rect 676 894 692 928
rect 626 884 692 894
rect 978 926 1044 936
rect 978 892 994 926
rect 1028 892 1044 926
rect 978 882 1044 892
rect 450 794 516 834
rect 1156 794 1228 834
rect 450 758 490 794
rect 1188 764 1228 794
rect 978 746 1044 756
rect 978 712 994 746
rect 1028 712 1044 746
rect 978 702 1044 712
rect 722 368 776 384
rect 722 334 732 368
rect 766 334 776 368
rect 722 318 776 334
rect 1074 326 1140 336
rect 1074 292 1090 326
rect 1124 292 1140 326
rect 1074 282 1140 292
rect 450 130 490 164
rect 450 90 516 130
rect 658 90 720 130
rect 680 60 720 90
rect 854 -174 908 -158
rect 854 -208 864 -174
rect 898 -208 908 -174
rect 854 -224 908 -208
rect 680 -272 720 -238
rect 1188 -272 1228 -238
rect 388 -416 412 -272
rect 1228 -416 1252 -272
<< viali >>
rect 414 1640 1200 1772
rect 538 1000 578 1600
rect 832 1000 930 1600
rect 1184 1000 1224 1600
rect 642 894 676 928
rect 994 892 1028 926
rect 450 164 490 758
rect 994 712 1028 746
rect 732 334 766 368
rect 1090 292 1124 326
rect 680 -238 720 60
rect 864 -208 898 -174
rect 1188 -238 1228 764
rect 412 -408 1228 -280
<< metal1 >>
rect 532 1778 584 1780
rect 348 1772 1260 1778
rect 348 1640 414 1772
rect 1200 1640 1260 1772
rect 348 1634 1260 1640
rect 532 1600 584 1634
rect 532 1000 538 1600
rect 578 1000 584 1600
rect 638 1580 684 1634
rect 826 1600 936 1634
rect 532 976 584 1000
rect 826 1000 832 1600
rect 930 1000 936 1600
rect 990 1578 1036 1634
rect 1178 1600 1230 1634
rect 616 934 692 938
rect 616 880 624 934
rect 684 880 692 934
rect 616 876 692 880
rect 726 936 772 980
rect 826 976 936 1000
rect 1178 1000 1184 1600
rect 1224 1000 1230 1600
rect 726 926 1044 936
rect 726 892 994 926
rect 1028 892 1044 926
rect 726 882 1044 892
rect 444 758 496 834
rect 444 164 450 758
rect 490 164 496 758
rect 726 756 772 882
rect 550 746 1044 756
rect 550 712 994 746
rect 1028 712 1044 746
rect 550 702 1044 712
rect 550 634 596 702
rect 726 634 772 702
rect 1078 634 1124 978
rect 1178 974 1230 1000
rect 1182 764 1234 834
rect 638 270 684 434
rect 718 378 780 384
rect 718 314 722 378
rect 776 314 780 378
rect 718 308 780 314
rect 814 280 860 434
rect 902 280 948 434
rect 990 280 1036 434
rect 1074 336 1150 340
rect 1074 282 1082 336
rect 1142 282 1150 336
rect 1074 278 1150 282
rect 638 224 814 270
rect 444 136 496 164
rect 444 84 726 136
rect 674 60 726 84
rect 674 -238 680 60
rect 720 -238 726 60
rect 850 -164 912 -158
rect 850 -228 854 -164
rect 908 -228 912 -164
rect 850 -234 912 -228
rect 674 -272 726 -238
rect 990 -272 1036 -120
rect 1182 -238 1188 764
rect 1228 -238 1234 764
rect 1182 -272 1234 -238
rect 348 -280 1260 -272
rect 348 -408 412 -280
rect 1228 -408 1260 -280
rect 348 -416 1260 -408
<< via1 >>
rect 624 928 684 934
rect 624 894 642 928
rect 642 894 676 928
rect 676 894 684 928
rect 624 880 684 894
rect 722 368 776 378
rect 722 334 732 368
rect 732 334 766 368
rect 766 334 776 368
rect 722 314 776 334
rect 1082 326 1142 336
rect 1082 292 1090 326
rect 1090 292 1124 326
rect 1124 292 1142 326
rect 1082 282 1142 292
rect 854 -174 908 -164
rect 854 -208 864 -174
rect 864 -208 898 -174
rect 898 -208 908 -174
rect 854 -228 908 -208
<< metal2 >>
rect 348 934 692 938
rect 348 880 624 934
rect 684 880 692 934
rect 348 876 692 880
rect 348 368 408 876
rect 718 378 780 384
rect 718 368 722 378
rect 348 314 722 368
rect 776 314 780 378
rect 348 308 780 314
rect 1074 336 1150 340
rect 1074 282 1082 336
rect 1142 282 1150 336
rect 1074 278 1150 282
rect 850 -164 912 -158
rect 850 -228 854 -164
rect 908 -228 912 -164
rect 850 -234 912 -228
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1730191042
transform 1 0 617 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1730191042
transform 1 0 705 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1730191042
transform 1 0 793 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1730191042
transform 1 0 881 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1730191042
transform 1 0 969 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1730191042
transform 1 0 1057 0 1 534
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_TC9PQS  sky130_fd_pr__nfet_01v8_TC9PQS_0
timestamp 1731171178
transform 1 0 881 0 1 80
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PQS  sky130_fd_pr__nfet_01v8_TC9PQS_1
timestamp 1731171178
transform 1 0 969 0 1 80
box -73 -226 73 226
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 705 0 1 1280
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_1
timestamp 1730191042
transform 1 0 1057 0 1 1278
box -109 -362 109 362
<< labels >>
rlabel metal2 348 732 400 784 0 in
port 1 nsew
rlabel metal2 850 -210 902 -158 0 t0
port 2 nsew
rlabel metal2 1074 288 1126 340 0 t1
port 3 nsew
rlabel metal1 348 1726 400 1778 0 VDD
port 5 nsew
rlabel metal1 348 -324 400 -272 0 VSS
port 6 nsew
rlabel metal1 1078 882 1124 928 0 out
port 4 nsew
<< end >>
