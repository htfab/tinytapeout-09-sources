magic
tech sky130A
magscale 1 2
timestamp 1730493024
<< error_p >>
rect -125 481 -67 487
rect 67 481 125 487
rect -125 447 -113 481
rect 67 447 79 481
rect -125 441 -67 447
rect 67 441 125 447
rect -221 -447 -163 -441
rect -29 -447 29 -441
rect 163 -447 221 -441
rect -221 -481 -209 -447
rect -29 -481 -17 -447
rect 163 -481 175 -447
rect -221 -487 -163 -481
rect -29 -487 29 -481
rect 163 -487 221 -481
<< nwell >>
rect -407 -619 407 619
<< pmos >>
rect -207 -400 -177 400
rect -111 -400 -81 400
rect -15 -400 15 400
rect 81 -400 111 400
rect 177 -400 207 400
<< pdiff >>
rect -269 388 -207 400
rect -269 -388 -257 388
rect -223 -388 -207 388
rect -269 -400 -207 -388
rect -177 388 -111 400
rect -177 -388 -161 388
rect -127 -388 -111 388
rect -177 -400 -111 -388
rect -81 388 -15 400
rect -81 -388 -65 388
rect -31 -388 -15 388
rect -81 -400 -15 -388
rect 15 388 81 400
rect 15 -388 31 388
rect 65 -388 81 388
rect 15 -400 81 -388
rect 111 388 177 400
rect 111 -388 127 388
rect 161 -388 177 388
rect 111 -400 177 -388
rect 207 388 269 400
rect 207 -388 223 388
rect 257 -388 269 388
rect 207 -400 269 -388
<< pdiffc >>
rect -257 -388 -223 388
rect -161 -388 -127 388
rect -65 -388 -31 388
rect 31 -388 65 388
rect 127 -388 161 388
rect 223 -388 257 388
<< nsubdiff >>
rect -371 549 -275 583
rect 275 549 371 583
rect -371 487 -337 549
rect 337 487 371 549
rect -371 -549 -337 -487
rect 337 -549 371 -487
rect -371 -583 -275 -549
rect 275 -583 371 -549
<< nsubdiffcont >>
rect -275 549 275 583
rect -371 -487 -337 487
rect 337 -487 371 487
rect -275 -583 275 -549
<< poly >>
rect -129 481 -63 497
rect -129 447 -113 481
rect -79 447 -63 481
rect -129 431 -63 447
rect 63 481 129 497
rect 63 447 79 481
rect 113 447 129 481
rect 63 431 129 447
rect -207 400 -177 426
rect -111 400 -81 431
rect -15 400 15 426
rect 81 400 111 431
rect 177 400 207 426
rect -207 -431 -177 -400
rect -111 -426 -81 -400
rect -15 -431 15 -400
rect 81 -426 111 -400
rect 177 -431 207 -400
rect -225 -447 -159 -431
rect -225 -481 -209 -447
rect -175 -481 -159 -447
rect -225 -497 -159 -481
rect -33 -447 33 -431
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect -33 -497 33 -481
rect 159 -447 225 -431
rect 159 -481 175 -447
rect 209 -481 225 -447
rect 159 -497 225 -481
<< polycont >>
rect -113 447 -79 481
rect 79 447 113 481
rect -209 -481 -175 -447
rect -17 -481 17 -447
rect 175 -481 209 -447
<< locali >>
rect -371 549 -275 583
rect 275 549 371 583
rect -371 487 -337 549
rect 337 487 371 549
rect -129 447 -113 481
rect -79 447 -63 481
rect 63 447 79 481
rect 113 447 129 481
rect -257 388 -223 404
rect -257 -404 -223 -388
rect -161 388 -127 404
rect -161 -404 -127 -388
rect -65 388 -31 404
rect -65 -404 -31 -388
rect 31 388 65 404
rect 31 -404 65 -388
rect 127 388 161 404
rect 127 -404 161 -388
rect 223 388 257 404
rect 223 -404 257 -388
rect -225 -481 -209 -447
rect -175 -481 -159 -447
rect -33 -481 -17 -447
rect 17 -481 33 -447
rect 159 -481 175 -447
rect 209 -481 225 -447
rect -371 -549 -337 -487
rect 337 -549 371 -487
rect -371 -583 -275 -549
rect 275 -583 371 -549
<< viali >>
rect -113 447 -79 481
rect 79 447 113 481
rect -257 -388 -223 388
rect -161 -388 -127 388
rect -65 -388 -31 388
rect 31 -388 65 388
rect 127 -388 161 388
rect 223 -388 257 388
rect -209 -481 -175 -447
rect -17 -481 17 -447
rect 175 -481 209 -447
<< metal1 >>
rect -125 481 -67 487
rect -125 447 -113 481
rect -79 447 -67 481
rect -125 441 -67 447
rect 67 481 125 487
rect 67 447 79 481
rect 113 447 125 481
rect 67 441 125 447
rect -263 388 -217 400
rect -263 -388 -257 388
rect -223 -388 -217 388
rect -263 -400 -217 -388
rect -167 388 -121 400
rect -167 -388 -161 388
rect -127 -388 -121 388
rect -167 -400 -121 -388
rect -71 388 -25 400
rect -71 -388 -65 388
rect -31 -388 -25 388
rect -71 -400 -25 -388
rect 25 388 71 400
rect 25 -388 31 388
rect 65 -388 71 388
rect 25 -400 71 -388
rect 121 388 167 400
rect 121 -388 127 388
rect 161 -388 167 388
rect 121 -400 167 -388
rect 217 388 263 400
rect 217 -388 223 388
rect 257 -388 263 388
rect 217 -400 263 -388
rect -221 -447 -163 -441
rect -221 -481 -209 -447
rect -175 -481 -163 -447
rect -221 -487 -163 -481
rect -29 -447 29 -441
rect -29 -481 -17 -447
rect 17 -481 29 -447
rect -29 -487 29 -481
rect 163 -447 221 -441
rect 163 -481 175 -447
rect 209 -481 221 -447
rect 163 -487 221 -481
<< properties >>
string FIXED_BBOX -354 -566 354 566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
