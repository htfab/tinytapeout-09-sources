magic
tech sky130A
magscale 1 2
timestamp 1728214159
<< error_p >>
rect -29 672 29 678
rect -29 638 -17 672
rect -29 632 29 638
rect -125 -638 -67 -632
rect 67 -638 125 -632
rect -125 -672 -113 -638
rect 67 -672 79 -638
rect -125 -678 -67 -672
rect 67 -678 125 -672
<< pwell >>
rect -311 -810 311 810
<< nmos >>
rect -111 -600 -81 600
rect -15 -600 15 600
rect 81 -600 111 600
<< ndiff >>
rect -173 588 -111 600
rect -173 -588 -161 588
rect -127 -588 -111 588
rect -173 -600 -111 -588
rect -81 588 -15 600
rect -81 -588 -65 588
rect -31 -588 -15 588
rect -81 -600 -15 -588
rect 15 588 81 600
rect 15 -588 31 588
rect 65 -588 81 588
rect 15 -600 81 -588
rect 111 588 173 600
rect 111 -588 127 588
rect 161 -588 173 588
rect 111 -600 173 -588
<< ndiffc >>
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
<< psubdiff >>
rect -275 740 -179 774
rect 179 740 275 774
rect -275 678 -241 740
rect 241 678 275 740
rect -275 -740 -241 -678
rect 241 -740 275 -678
rect -275 -774 -179 -740
rect 179 -774 275 -740
<< psubdiffcont >>
rect -179 740 179 774
rect -275 -678 -241 678
rect 241 -678 275 678
rect -179 -774 179 -740
<< poly >>
rect -33 672 33 688
rect -33 638 -17 672
rect 17 638 33 672
rect -111 600 -81 626
rect -33 622 33 638
rect -15 600 15 622
rect 81 600 111 626
rect -111 -622 -81 -600
rect -129 -638 -63 -622
rect -15 -626 15 -600
rect 81 -622 111 -600
rect -129 -672 -113 -638
rect -79 -672 -63 -638
rect -129 -688 -63 -672
rect 63 -638 129 -622
rect 63 -672 79 -638
rect 113 -672 129 -638
rect 63 -688 129 -672
<< polycont >>
rect -17 638 17 672
rect -113 -672 -79 -638
rect 79 -672 113 -638
<< locali >>
rect -275 740 -179 774
rect 179 740 275 774
rect -275 678 -241 740
rect 241 678 275 740
rect -33 638 -17 672
rect 17 638 33 672
rect -161 588 -127 604
rect -161 -604 -127 -588
rect -65 588 -31 604
rect -65 -604 -31 -588
rect 31 588 65 604
rect 31 -604 65 -588
rect 127 588 161 604
rect 127 -604 161 -588
rect -129 -672 -113 -638
rect -79 -672 -63 -638
rect 63 -672 79 -638
rect 113 -672 129 -638
rect -275 -740 -241 -678
rect 241 -740 275 -678
rect -275 -774 -179 -740
rect 179 -774 275 -740
<< viali >>
rect -17 638 17 672
rect -161 -588 -127 588
rect -65 -588 -31 588
rect 31 -588 65 588
rect 127 -588 161 588
rect -113 -672 -79 -638
rect 79 -672 113 -638
<< metal1 >>
rect -29 672 29 678
rect -29 638 -17 672
rect 17 638 29 672
rect -29 632 29 638
rect -167 588 -121 600
rect -167 -588 -161 588
rect -127 -588 -121 588
rect -167 -600 -121 -588
rect -71 588 -25 600
rect -71 -588 -65 588
rect -31 -588 -25 588
rect -71 -600 -25 -588
rect 25 588 71 600
rect 25 -588 31 588
rect 65 -588 71 588
rect 25 -600 71 -588
rect 121 588 167 600
rect 121 -588 127 588
rect 161 -588 167 588
rect 121 -600 167 -588
rect -125 -638 -67 -632
rect -125 -672 -113 -638
rect -79 -672 -67 -638
rect -125 -678 -67 -672
rect 67 -638 125 -632
rect 67 -672 79 -638
rect 113 -672 125 -638
rect 67 -678 125 -672
<< properties >>
string FIXED_BBOX -258 -757 258 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
