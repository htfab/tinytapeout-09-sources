magic
tech sky130A
magscale 1 2
timestamp 1730821126
<< nwell >>
rect -444 1084 836 1380
rect -444 360 -292 1084
rect 190 1080 378 1084
rect 190 970 268 1080
rect 270 1064 378 1080
rect 474 1064 538 1084
rect -198 360 -80 396
rect -22 360 96 396
rect 188 388 268 970
rect 190 360 268 388
rect 284 360 378 1064
rect 384 360 458 396
rect 718 360 836 1084
<< pwell >>
rect -444 -142 836 360
<< psubdiff >>
rect -348 272 -310 296
rect -348 -46 -310 -10
rect 208 272 246 296
rect 208 -46 246 -10
rect 764 272 802 296
rect 764 -46 802 -10
rect -382 -142 -358 -46
rect 812 -142 836 -46
<< nsubdiff >>
rect -346 1248 -322 1344
rect 768 1248 800 1344
rect -346 1214 -310 1248
rect -346 418 -310 442
rect 208 1214 246 1248
rect 208 418 246 442
rect 764 1214 800 1248
rect 764 418 800 442
<< psubdiffcont >>
rect -348 -10 -310 272
rect 208 -10 246 272
rect 764 -10 802 272
rect -358 -142 812 -46
<< nsubdiffcont >>
rect -322 1248 768 1344
rect -346 442 -310 1214
rect 208 442 246 1214
rect 764 442 800 1214
<< poly >>
rect -198 386 -168 396
rect -110 386 -80 396
rect -198 374 -80 386
rect -198 338 -158 374
rect -122 338 -80 374
rect -198 326 -80 338
rect -198 318 -168 326
rect -110 318 -80 326
rect -22 386 8 396
rect 66 386 96 396
rect -22 374 96 386
rect -22 338 18 374
rect 54 338 96 374
rect -22 326 96 338
rect -22 318 8 326
rect 66 318 96 326
rect 358 386 388 396
rect 446 386 476 396
rect 358 374 476 386
rect 358 338 398 374
rect 434 338 476 374
rect 358 326 476 338
rect 358 318 388 326
rect 446 318 476 326
rect 534 386 564 396
rect 622 386 652 396
rect 534 374 652 386
rect 534 338 576 374
rect 612 338 652 374
rect 534 326 652 338
rect 534 318 564 326
rect 622 318 652 326
<< polycont >>
rect -158 338 -122 374
rect 18 338 54 374
rect 398 338 434 374
rect 576 338 612 374
<< locali >>
rect -346 1248 -322 1344
rect 768 1248 800 1344
rect -346 1214 -310 1248
rect -346 418 -310 442
rect 208 1214 246 1248
rect 208 418 246 442
rect 764 1214 800 1248
rect 764 418 800 442
rect -174 338 -158 374
rect -122 338 -106 374
rect 2 338 18 374
rect 54 338 70 374
rect 382 338 398 374
rect 434 338 450 374
rect 560 338 576 374
rect 612 338 628 374
rect -348 272 -310 296
rect -348 -46 -310 -10
rect 208 272 246 296
rect 208 -46 246 -10
rect 764 272 802 296
rect 764 -46 802 -10
rect -382 -142 -358 -46
rect 812 -142 836 -46
<< viali >>
rect -322 1254 768 1338
rect -346 442 -310 1214
rect 764 442 800 1214
rect -158 338 -122 374
rect 18 338 54 374
rect 398 338 434 374
rect 576 338 612 374
rect -348 -10 -310 272
rect 764 -10 802 272
rect -358 -136 812 -52
<< metal1 >>
rect -444 1338 836 1344
rect -444 1254 -322 1338
rect 768 1254 836 1338
rect -444 1248 836 1254
rect -352 1214 -304 1248
rect -352 442 -346 1214
rect -310 442 -304 1214
rect -268 1214 -204 1220
rect -268 1162 -262 1214
rect -210 1162 -204 1214
rect -268 1156 -204 1162
rect -250 1022 -204 1156
rect -162 1022 -116 1248
rect -82 1122 -18 1128
rect -82 1070 -76 1122
rect -24 1070 -18 1122
rect -82 1064 -18 1070
rect -74 1022 -28 1064
rect 14 1022 60 1248
rect 188 1214 252 1220
rect 188 1162 194 1214
rect 246 1162 252 1214
rect 92 1122 156 1128
rect 92 1070 98 1122
rect 150 1070 156 1122
rect 92 1064 156 1070
rect 102 1022 148 1064
rect 188 964 252 1162
rect 394 1022 440 1248
rect 570 1022 616 1248
rect 758 1214 806 1248
rect 188 912 194 964
rect 246 912 252 964
rect 188 906 252 912
rect 208 442 246 906
rect 758 442 764 1214
rect 800 442 806 1214
rect -352 418 -304 442
rect -354 272 -304 296
rect -250 292 -204 422
rect -172 382 -108 386
rect -172 330 -166 382
rect -114 330 -108 382
rect -172 326 -108 330
rect -74 292 -28 422
rect 4 382 68 386
rect 4 330 10 382
rect 62 330 68 382
rect 4 326 68 330
rect 102 292 148 422
rect 306 292 352 422
rect 384 382 448 386
rect 384 330 390 382
rect 442 330 448 382
rect 384 326 448 330
rect 482 292 528 422
rect 562 382 626 386
rect 562 330 568 382
rect 620 330 626 382
rect 562 326 626 330
rect 658 292 704 422
rect 758 418 806 442
rect -354 -10 -348 272
rect -310 -10 -304 272
rect 758 272 808 296
rect -354 -46 -304 -10
rect -162 -46 -116 94
rect 14 -46 60 92
rect 102 88 148 92
rect 306 50 352 92
rect 102 44 352 50
rect 102 -8 108 44
rect 160 4 352 44
rect 160 -8 166 4
rect 102 -14 166 -8
rect 394 -46 440 92
rect 482 50 528 92
rect 474 44 538 50
rect 474 -8 480 44
rect 532 -8 538 44
rect 474 -14 538 -8
rect 570 -46 616 92
rect 658 50 704 92
rect 658 44 722 50
rect 658 -8 664 44
rect 716 -8 722 44
rect 658 -14 722 -8
rect 758 -10 764 272
rect 802 -10 808 272
rect 758 -46 808 -10
rect -444 -52 836 -46
rect -444 -136 -358 -52
rect 812 -136 836 -52
rect -444 -142 836 -136
<< via1 >>
rect -262 1162 -210 1214
rect -76 1070 -24 1122
rect 194 1162 246 1214
rect 98 1070 150 1122
rect 194 912 246 964
rect -166 374 -114 382
rect -166 338 -158 374
rect -158 338 -122 374
rect -122 338 -114 374
rect -166 330 -114 338
rect 10 374 62 382
rect 10 338 18 374
rect 18 338 54 374
rect 54 338 62 374
rect 10 330 62 338
rect 390 374 442 382
rect 390 338 398 374
rect 398 338 434 374
rect 434 338 442 374
rect 390 330 442 338
rect 568 374 620 382
rect 568 338 576 374
rect 576 338 612 374
rect 612 338 620 374
rect 568 330 620 338
rect 108 -8 160 44
rect 480 -8 532 44
rect 664 -8 716 44
<< metal2 >>
rect -444 1214 252 1220
rect -444 1162 -262 1214
rect -210 1162 194 1214
rect 246 1162 252 1214
rect -444 1156 252 1162
rect 474 1156 836 1220
rect 474 1128 538 1156
rect -82 1122 538 1128
rect -82 1070 -76 1122
rect -24 1070 98 1122
rect 150 1070 538 1122
rect -82 1064 538 1070
rect 188 964 252 970
rect 188 912 194 964
rect 246 912 252 964
rect 188 388 252 912
rect -444 382 96 388
rect -444 330 -166 382
rect -114 330 10 382
rect 62 330 96 382
rect -444 324 96 330
rect 188 382 654 388
rect 188 330 390 382
rect 442 330 568 382
rect 620 330 654 382
rect 188 324 654 330
rect -444 50 -380 324
rect -444 44 166 50
rect -444 -8 108 44
rect 160 -8 166 44
rect -444 -14 166 -8
rect 474 44 836 50
rect 474 -8 480 44
rect 532 -8 664 44
rect 716 -8 836 44
rect 474 -14 836 -8
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1730191042
transform 1 0 81 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1730191042
transform 1 0 -7 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1730191042
transform 1 0 -95 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1730191042
transform 1 0 -183 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_4
timestamp 1730191042
transform 1 0 373 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_5
timestamp 1730191042
transform 1 0 461 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_6
timestamp 1730191042
transform 1 0 549 0 1 192
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_7
timestamp 1730191042
transform 1 0 637 0 1 192
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_0
timestamp 1730191042
transform 1 0 81 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_1
timestamp 1730191042
transform 1 0 -7 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_2
timestamp 1730191042
transform 1 0 -95 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_3
timestamp 1730191042
transform 1 0 -183 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_4
timestamp 1730191042
transform 1 0 461 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_5
timestamp 1730191042
transform 1 0 373 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_6
timestamp 1730191042
transform 1 0 637 0 1 722
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_2K9SAN  sky130_fd_pr__pfet_01v8_2K9SAN_7
timestamp 1730191042
transform 1 0 549 0 1 722
box -109 -362 109 362
<< labels >>
rlabel metal2 -444 -14 -380 50 0 in_2
port 2 nsew
rlabel metal2 772 -14 836 50 0 out_2
port 4 nsew
rlabel metal2 -382 1156 -318 1220 0 in_1
port 1 nsew
rlabel nwell -382 1280 -318 1344 0 VDD
port 5 nsew
rlabel metal1 -442 -110 -378 -46 0 VSS
port 6 nsew
rlabel metal2 772 1156 836 1220 0 out_1
port 3 nsew
<< end >>
