magic
tech sky130A
magscale 1 2
timestamp 1730911581
<< nwell >>
rect 2751 840 4479 1299
rect 2642 802 4479 840
rect 2642 -399 2852 802
<< pwell >>
rect 5119 -871 5255 -699
<< locali >>
rect 542 1679 5837 1713
rect 542 1617 566 1679
rect 539 1610 566 1617
rect 5778 1610 5837 1679
rect 539 1573 2799 1610
rect 539 1522 1386 1573
rect 2752 817 2799 1573
rect 3029 1573 5837 1610
rect 3029 817 3088 1573
rect 2752 778 3088 817
rect 5029 -1230 5544 -1031
rect 547 -1267 5863 -1230
rect 547 -1374 586 -1267
rect 5836 -1374 5863 -1267
rect 547 -1403 5863 -1374
<< viali >>
rect 566 1610 5778 1679
rect 2799 817 3029 1610
rect 586 -1374 5836 -1267
<< metal1 >>
rect 542 1679 5837 1713
rect 542 1610 566 1679
rect 5778 1610 5837 1679
rect 542 1573 2799 1610
rect 736 1421 1118 1573
rect 1536 1465 1913 1507
rect 2225 1465 2602 1507
rect 645 733 688 1381
rect 1164 733 1207 1376
rect 645 370 1207 733
rect 645 -114 688 370
rect 570 -187 688 -114
rect 867 -93 919 -87
rect 867 -151 919 -145
rect 1164 -150 1207 370
rect 1430 -81 1518 1403
rect 1622 76 1800 1465
rect 1944 1397 2007 1399
rect 878 -183 908 -151
rect 570 -1228 669 -187
rect 873 -219 914 -183
rect 1206 -192 1207 -150
rect 1374 -169 1518 -81
rect 1608 -124 1811 76
rect 1944 -93 2193 1397
rect 2317 448 2495 1465
rect 2316 124 2496 448
rect 2317 42 2495 124
rect 740 -248 1118 -219
rect 1374 -616 1448 -169
rect 1622 -226 1800 -124
rect 1944 -145 2043 -93
rect 2095 -145 2193 -93
rect 1944 -163 2193 -145
rect 2302 -158 2508 42
rect 2634 -154 2697 1403
rect 2752 817 2799 1573
rect 3029 1573 5837 1610
rect 3029 1326 3088 1573
rect 3255 1326 4240 1328
rect 3029 1230 4240 1326
rect 3029 817 3088 1230
rect 3156 1105 3207 1113
rect 3255 1106 4240 1230
rect 3150 1050 3156 1105
rect 3211 1050 3217 1105
rect 3156 1047 3207 1050
rect 3261 1010 4232 1050
rect 4294 1047 4345 1113
rect 2752 778 3088 817
rect 3261 701 3790 706
rect 3007 698 3790 701
rect 3001 666 3790 698
rect 3007 665 3790 666
rect 2764 588 2770 643
rect 2825 588 2831 643
rect 1944 -167 2007 -163
rect 2316 -186 2498 -158
rect 2634 -163 2700 -154
rect 1539 -268 1916 -226
rect 2314 -227 2516 -186
rect 2225 -269 2602 -227
rect 2661 -615 2700 -163
rect 2778 -513 2816 588
rect 2902 342 2976 609
rect 3247 342 3516 665
rect 3893 599 3991 1010
rect 4105 701 4232 706
rect 4105 665 4871 701
rect 2902 65 3516 342
rect 2902 -81 2976 65
rect 2901 -180 2976 -81
rect 2778 -551 2841 -513
rect 854 -647 1618 -616
rect 1934 -647 2700 -615
rect 792 -776 826 -698
rect 1082 -776 1240 -647
rect 792 -821 1240 -776
rect 792 -837 1026 -821
rect 775 -840 1026 -837
rect 758 -873 1026 -840
rect 1078 -873 1240 -821
rect 758 -1009 1240 -873
rect 758 -1075 826 -1009
rect 758 -1084 803 -1075
rect 1082 -1123 1240 -1009
rect 1656 -1068 1907 -703
rect 2215 -730 2483 -647
rect 2803 -653 2841 -551
rect 2215 -968 2765 -730
rect 2215 -1027 2517 -968
rect 2576 -1027 2765 -968
rect 2215 -1049 2765 -1027
rect 855 -1154 1619 -1123
rect 758 -1228 803 -1226
rect 1738 -1228 1836 -1068
rect 2215 -1125 2483 -1049
rect 2806 -1122 2841 -653
rect 2901 -697 2960 -180
rect 3247 -229 3516 65
rect 3807 -166 4061 599
rect 4357 -229 4626 665
rect 5061 606 5156 1573
rect 5421 1412 5557 1573
rect 5641 1468 5708 1518
rect 5421 1312 5641 1412
rect 5235 668 5302 718
rect 4907 604 4975 605
rect 4897 -174 4975 604
rect 5061 457 5231 606
rect 5128 -166 5231 457
rect 5296 -95 5391 616
rect 5296 -169 5428 -95
rect 5528 -159 5641 1312
rect 5704 -57 5849 1407
rect 5704 -163 5864 -57
rect 3008 -261 4872 -229
rect 4907 -547 4975 -174
rect 5237 -547 5321 -218
rect 4907 -578 5321 -547
rect 4922 -601 5321 -578
rect 3030 -649 3798 -613
rect 4109 -649 4877 -613
rect 2901 -838 2997 -697
rect 2915 -1074 2997 -838
rect 3290 -968 3481 -649
rect 3290 -1027 3347 -968
rect 3406 -1027 3481 -968
rect 1941 -1157 2707 -1125
rect 2803 -1228 2841 -1122
rect 3290 -1128 3481 -1027
rect 3823 -1073 4082 -699
rect 4379 -821 4570 -649
rect 4922 -685 4975 -601
rect 5237 -656 5321 -601
rect 5368 -408 5428 -169
rect 5627 -314 5730 -216
rect 5627 -407 5729 -314
rect 5790 -320 5864 -163
rect 5554 -408 5729 -407
rect 5368 -489 5729 -408
rect 5368 -657 5428 -489
rect 5554 -492 5729 -489
rect 5627 -514 5729 -492
rect 5627 -654 5730 -514
rect 5775 -520 5975 -320
rect 4379 -873 4450 -821
rect 4502 -873 4570 -821
rect 3020 -1164 3788 -1128
rect 3897 -1228 4008 -1073
rect 4379 -1123 4570 -873
rect 4907 -1075 4975 -685
rect 5380 -694 5428 -657
rect 5119 -833 5255 -699
rect 5117 -871 5255 -833
rect 5315 -760 5428 -694
rect 5790 -697 5864 -520
rect 5315 -871 5405 -760
rect 5117 -1031 5188 -871
rect 5253 -972 5320 -922
rect 5577 -926 5657 -705
rect 5513 -1031 5657 -926
rect 5029 -1067 5657 -1031
rect 5714 -762 5864 -697
rect 4109 -1159 4877 -1123
rect 5029 -1155 5590 -1067
rect 5714 -1070 5863 -762
rect 5029 -1228 5522 -1155
rect 5656 -1170 5723 -1120
rect 547 -1267 5868 -1228
rect 547 -1374 586 -1267
rect 5836 -1374 5868 -1267
rect 547 -1403 5868 -1374
<< via1 >>
rect 867 -145 919 -93
rect 2043 -145 2095 -93
rect 3156 1050 3211 1105
rect 2770 588 2825 643
rect 1026 -873 1078 -821
rect 2517 -1027 2576 -968
rect 3347 -1027 3406 -968
rect 4450 -873 4502 -821
<< metal2 >>
rect 3156 1105 3211 1111
rect 2770 1050 3156 1105
rect 2770 643 2825 1050
rect 3156 1044 3211 1050
rect 2770 582 2825 588
rect 861 -145 867 -93
rect 919 -104 925 -93
rect 2037 -104 2043 -93
rect 919 -134 2043 -104
rect 919 -145 925 -134
rect 2037 -145 2043 -134
rect 2095 -145 2101 -93
rect 1020 -873 1026 -821
rect 1078 -826 1084 -821
rect 4444 -826 4450 -821
rect 1078 -868 4450 -826
rect 1078 -873 1084 -868
rect 4444 -873 4450 -868
rect 4502 -873 4508 -821
rect 2511 -1027 2517 -968
rect 2576 -1027 3347 -968
rect 3406 -1027 3412 -968
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM1
timestamp 1730892491
transform 1 0 1238 0 1 -886
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM2
timestamp 1730892491
transform 1 0 2324 0 1 -886
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM3
timestamp 1730892491
transform 1 0 3410 0 1 -886
box -596 -410 596 410
use sky130_fd_pr__nfet_01v8_lvt_FMZK9W  XM4
timestamp 1730892491
transform 1 0 4496 0 1 -886
box -596 -410 596 410
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM5
timestamp 1730892491
transform 1 0 1730 0 1 619
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_GWPMZG  XM6
timestamp 1730892491
transform 1 0 2416 0 1 619
box -396 -1019 396 1019
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM7
timestamp 1730892491
transform 1 0 3392 0 1 218
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_GGY9VD  XM8
timestamp 1730892491
transform 0 1 929 -1 0 596
box -996 -419 996 419
use sky130_fd_pr__pfet_01v8_lvt_ZQZ9VD  XM9
timestamp 1730892491
transform 1 0 4478 0 1 218
box -596 -619 596 619
use sky130_fd_pr__pfet_01v8_UGSVTG  XM10
timestamp 1730892491
transform 0 1 3752 -1 0 1079
box -211 -719 211 719
use sky130_fd_pr__pfet_01v8_XGASDL#0  XM11
timestamp 1730892491
transform 1 0 5268 0 1 221
box -211 -619 211 619
use sky130_fd_pr__nfet_01v8_648S5X#0  XM12
timestamp 1730892491
transform 1 0 5285 0 1 -785
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_UGACMG  XM13
timestamp 1730909037
transform 1 0 5673 0 1 622
box -211 -1019 211 1019
use sky130_fd_pr__nfet_01v8_ATLS57#0  XM14
timestamp 1730892491
transform 1 0 5690 0 1 -884
box -211 -410 211 410
<< labels >>
flabel metal1 5775 -520 5975 -320 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 5201 -1347 5401 -1147 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 2801 1463 3001 1663 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1611 -124 1811 76 0 FreeSans 256 0 0 0 in+
port 3 nsew
flabel metal1 2308 -158 2508 42 0 FreeSans 256 0 0 0 in-
port 4 nsew
<< end >>
